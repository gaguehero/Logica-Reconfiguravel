`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FRCRL+bzJpjrhpVLeYuwbH+fQ7cNyz7dW5pr/v860XGpwXN9jueTGVlRjaUB6XSn
uVE1/03O9dsORn1+RzjUamZ41a3nqVdNTMnjHG4fU28HPN12ct1THHSZYIpGfUGC
ISoVAaj+rTKCbA/C+YFA4uJnfb7sh1NKTOWAMZeHwtGYPCwpbggsERPWWtZ6/HUn
Wa9rvxYAIu9DDczkcQIHlZ44EmWboUBopWJUn86cx4a2Qz8JQpkfXHf9HFiDlsAV
8NEjobFpjJp1IPLmxkre7k2pDgVVCzavI+V9v05sHUiKWdqC8F9AfInWHzqL9EFt
vdghrF0dexiXMEon1NYuIlSNfnAjueMIwSJIpqknxYZK2UYHR1dyJf/D9yvwC3DA
fg2rmbEYKEzV6ixZ+HFB2oXwUuKHPh4NMHkQ4xslNIOWxe+j5uqMY6UeXLpc8fla
TPg/Pw+tQKCtEgEvrvBqj4OIDcbV+e258kv32TN0Asq2FU8iY1vhf21vkd5I+2/k
tQ/v6EJ4Vtp4Xb79pSiHnx0efQvNv5r38Ng/rNEPugKz310Ns8CvO58kVc8c4t6t
+/wVBOc+lDokB89RNZLrbMaXOI+BSk+dKlTMZ2gYBVvDOhLQvw4Jb4wGg/bK1OhJ
wuQxfXl8cWPLfb7Y6iiNyLLeI/EPwpVpAq+K66p52V+tAmQyfcyeWy9F8m15xGsz
lxCgqQ1Ce9Yqk/7zR6vioqdmAP9OxKzOToNSHK03crM=
`protect END_PROTECTED
