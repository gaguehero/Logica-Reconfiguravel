`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r84n81xy5Zi2gAL2iCTtMM0F8Mww3JRc206UsNHeQl834IQx2IHrD2hAdurvzALL
aiiCE4h99mgoDw2Kfi8/mdEpZYJH62YImgDlZ65dRZD3ax8DMVQKVdI2lv4DTFBA
aH57fyovXDt/nm6JfTINaz60pHDQvzHCP04Q+Ax0W/JgbS5sdPWevtFxPGdL+36+
xhhkq10aSj7ywJacrkLBKcVjdxNJSUT0XC9aqWAvsfJ5tK1UHUzoF+b6pHf06PMZ
o195NCvlFZi/WZl0IUpdG/dKBHozxUG5uzvXxEESal5MzCigLPbNPUAW8txLwqVm
CJGtKW7fv5tqhcoRJisQxzLYjy/mDHvE1P4963JESSFTQKB+rYTUdTV2I8kMRWcv
sMPgQXjq/RbqnEJRDrH+4BF9GcB8ELY00xH011MsxOq3Iwyeh30JZhbqisF56wxj
ocfSNMHAUGDssBBG8ckqg54LFZpp/hpiyv+ALOEz9WfrFXb//AGAvc7mRk5ng/+x
oUMAwe65qDqpp6Sikug0XHmmwDyJEuXgcvU2uUJbhNvW2oLre8do3hJ4YndjQSsO
vrkhseLW9yNVtOXoI5gy981FzmvBiGzUYueiefrULP4GRDVfUxvsQn26jfZ+m/PG
585+HNrJ3xO7qhh5OBW35PKh4MB6Yd7fZGwaJ0HYVS7Q7MvKCn67OmDhjmb1SCPa
M4t+fLupd0RJdcd8iSzU1E4s4XT5ecyn7f5oomb7763eUlREIDNZW1u8HMatW6Gw
xTQN3a5ODeNeArlXUvJkvSMSPA8DNf46jwhxxo1fmmJvjA5u6TOLkMFl1+uGHWlu
9jnsag7P2IbzTHKMpW9HJXCEKkt+T59vPd36h8R4xp5dwTx2fddkCci+/UvRm2xp
fLGj45UzjZGIjuSWlXE/B/xoPPaeaaAsxdpINCkUajxnYe12uvOfZonHZQ0XfDA9
pSpcOkvpum+zBSq6sKt/cxB7RM4ce51duf2iw1t6jbrsZySfhOmrkj8VbnnnfQob
4GcsFuChvZ0fRGabEkC7DfJQ0dv4DZYO4dwgipjJvlGMwCT++ZBQ0Zxi36m6zFAJ
m3nijT+nwIG4HhbNtw4SAN7tMbbL8nzwRWIGoG4jY58vY5SoEcATmFKsHaLcYHmg
Vijw9H/6K3GtNwwfjuFIiNCin+niHz3EhKdLvhQyE5bj/5xjGvrBG/dmvL6QpZjG
pHL0+x2nyoBki6nMP6CKMcsc+Tk8hY4+ThveUIi43mI=
`protect END_PROTECTED
