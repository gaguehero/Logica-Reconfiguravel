`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31uwySNkMf309TUryLptDJhNqPxVmVbFoqDCLnq5YLp0Qx5PuPTcMbQ3ZYGFnTUq
wsRoiR4RNgk0jiKVBAAWrwbEH06WVPCcsieEXGzFBEuCAk46h2teOaf5Ipy9kwJf
iDu89OBvoGcdGZeu4uWATLz44DZI78zPbCdJIvC9KdqJyLHaNQ7hlh+/YY0Qn1QF
GGwmFi8ZYUXWVXD3WDDETEoUpURDk1Ly2V3fHJw17GsiwkpPIkAJo/nNoPxG3kNP
URRBC7KJtb9N9oLnVwOd7/J+w1KzpyLn+qzCiRxgqz4jZrjFHprlC3RHe5poTZtW
eB5IegSg7G2f2nXuhrdilxvcyGQx9FilFCqJnWfEDZw4FHfpkQb+OhnRMKRJLsFR
+lolXmxMOJAY6l/KNJwTFUGZMjrr0xWZVOlsvIi48aq0uMz1otSPpsRA0Mz2fDNw
nzv717sxMSb4B4qDs393RIIMxpDpQ9/8uOPLc1PLVkokFLWG7kMb5GOhVcnowz04
rsjaFDt9HIcW+IfyigdzGhy/kffkcT76KS6qtpW4SJVJZQPi14JoXclaqOiTBDTz
Rw6qSArGGiHBMn7tFYjU55gLvYdGZpVLXNGhmbfXKaj2hSC27frmuhdBJVwluIwa
piZKzyS9UU4daHV5cLwlowGia8kOPIlFNatJmY3Hp8x7E+CT6I2wALTCGLTKwHL0
jjifORo/yRmVbZMqckbv8rx4tC0MvdZaNcdx4UYvIR+Hvzzoop0Hpc/kVvRXlQWZ
BJWw42r0aSRrmSgWJXdAu9YhU0N2PIhwat5E3+k5i8I8wQXIFi4gEk8LwwqJ3tU+
XFHrkUlo7ku2ymT9iOdgi80SYUNnCfTzNa+wOKlsNLYuZ4x7PaVEsjig8L4s96+4
sRnRVGTzyw4hN76KqWhbAossnr0zY5JdEpVIN/Jnn5Bs/HHxIMwaJl1h3Nfxy0TD
t+7R7moBn/KzU4fighbkpeS8iO2sKnLZIXVkznoWIz39w1KzTrr28zvhADGO8y+p
mZn+h3TtxDusq0MstScnlCtShzmE5m7gcao23KmgyiYmcN9b0cXKtNfsa01pCiAn
gwbboE+jvjHAp+wicr7jKcpeN6q72X68AlyNC2Ixnm+ViWWhxRg/6L/GiyXbKeSm
ZRXlG51/ZMur0ZqK77LrBG47j6ScTuAusH3TOwo9RqMzy7SPgzGJYSn+zHDvD/6G
Vb//qnmM6ruyj46v4AC2v1/ivGZ/rNmh+MFzf/mOl8HZ6TFNPtCRykifWCbi1sbU
1A2QTIr4DS2CiBI3MAkfEtztmN+lsddczQqx6ZsjSEp2A/nAGInCSqjZWddaZtMN
xZADiiv4braQpMZumx/ya3xsEiS717a5Cg0qN5P2CxvvSp/NMccdx9ih2UIxmkOt
0OqYK47dMHm0OkrPA7LN1HpMkSIa+FY/BGuDko6LBN9lZfXiFgvpY47WuZysSIa5
xRZ91b6a3IuDYfEvC3ezU+vgwVH1TzU2Ng2XjR4Rsn/xfHWfHC1xOhu9izfjiBvk
B9sWFrbCRXZUZtF0mw+ATYjv7gmI9L7NLqPpNqeJiCT+CYKwRKZoZ3KsWrsW52Xz
u9bVPw2b3Sq7tLzsGCMsXzkm8uGMKPRl35dxbZ82x5dB/0DYECWkazUPGDisPFp7
kEdIk9WwoqG3hFC1njk2WSV/9JE0q8S1EMmb0nqObErAaD+V0g9sWEKDva+bQEmb
wsKwwOhXM6Wnm4CU1VHuhXMLiM4to8k5iR88Z/p4AkDQhapuHPu2vJX88o8qRIbF
Tey4hg7jbb3BRt4cKwEp9lsH8hOuBkcWeTmX1D7//h5xq+ogjOKHCbmbHqh73yas
WqQnZBPZyhsCZa2VEyn+JpYeQ4kawgbjPIpusNfRrNE/uMcdgEUWBXNTX6rY3Kl4
jKMKsXcNWeabyjm7lrjVzkitlJH5wU2Mvp8Iq98G5qsYttePRZvIZXZepXvj9e6f
3UEOD24IGmjOfujwaMd0jA==
`protect END_PROTECTED
