`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3aX2mXQfcj1mB4R9JIyOq6KBMKQLGht2LVlSu5hsk5SiMR0aCpkERtq+rEY3jXUO
g3K7y2oLRBj3w76GSuXjdYNTt2hSchHe4y9HeIWrQR1nzojxhZsAMVbN3wAL6lTS
H7Y5yBdl73q7tK3t7lCAbW+gO3XpU0sTznGpnXiCtZIUdwNOA9WjNJr4fAsN5g/D
1fWGJVV8GikJ4gZj/YtJQ3wqSoVwjMJaYgslpyDAlWwog/KdYJopQjUsG1c3AC5V
RUEsoHhwWVN/EfxaPfa97Xi12HbHYx7x5/UW+ixl6aduezPHQ4fKijmvUGHlMhig
U0RKEyEXJWnCghqz+v9+xQOEpTb+KqaO3uEoAcF8BpyEEL2EDhoTskHdW1I+QG3X
KLQaoHXFI7CT+NzB9+gvgVrvbGXzUCnYAYNlTMTW7n8hhUxzWkFxrhj8kT6KUyhm
AXytS7+umkIWh5jAUUSYDiolyErBzcrXyZRWik3SNUQ3hxnNRULZuqBparmxoAEk
goj+xXlmyUp30/2oL9TZqDuKh5VamCBXJfgwWbANjtVRm9RiGBFe6/I5oBcWb2Vj
iighWVoXsNdS+WxRWlhjbE4TSLt6zCSmN7eB3aXZsT8=
`protect END_PROTECTED
