`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9b6wkPJOOSGqiVVERX0Gx3slX4VZfETaQl1cwtqeV0LGS9Iw65FYyF5Z6Fw0khSn
44amVxoGyUMITiaDP5ILXgUGxiiRBopljG9itYFBmK9YwZrlKmzwOl0SWAHn3y8g
Wali4T2l9eI6m4MBOWlpkyVfY2iBTg1F1M8UlPNd5o3kQAMnPDHL6g4hHQMn9VwD
JjrdV7iXqLes6xkLg+lvP4HvJDAIGRcjC9S7KJL4B+eNAvfn06Ze3LFykZj3bBXt
JEzvLEkgH8hWNFwCndpwGpqr+P9d21OoiT8wuUqFPcJt+oQpiu5qp0KHPT4YVFXR
Uc1SS5JF2lWEcFSHqe31dX6iVvhjhcI9gX9vpn9bja/Uvy1QNfTqQJp4rTeU0vLY
CX2+CFwei/HbCVUitrh/3RBU0mO+stjvxbAm3vx+nPQe6U4I/k5jhmEIYGsG4lRV
i0z+Uez/941hPHJVfPy6GSugq5w52a13+RhKVv3eOmyMEYMIvJzBHjjZaq2u4hPQ
2H8src+/1Meb5iq5mDTRw79aKex0V9O6yDwzLeZufdP91LTwnibYPgy0kDzmDEk+
duh6Us5/946nk6p2MjRzbR9ve5rkWwWHJ8sBGXTWev9rTlyGbFzi/GTyir1JiZvT
1tNq8U9WzjKo5UgZPN5yMO6BHaf+XcpyKFO20MtdDqTxHEVizx0UnGxxS/i0xnYQ
+XQLGERSOga7oHdk7CaOU8F+lVz4jx6TOeWFHgTu/6IrClxtvTNzjrx6bfpYwAXn
ioLDEpExCHztZy32Dh1SO1Cs04mBsnsDOQMZhTMjN++1rfejaSgjFqScTGLvdYny
bIOxqKqVN4zaqQS/i1E1gmxAnbeaJYfvpSPsc5tV2U94+jFnZg6bKHe/1orDy70S
3tBY2a0BesrF2oS6VLWDWg5EUQpib5Lqla7vOGNfHKwTYZzNDvVOGM+RrOdqdTjz
nYMlILfVN7pHQL3Jeu2iJwbXKilstTDXiM1xv7WYDVjYXYdHcLHKouVVh9PpenMY
ZtJNH5z/Zf4V2kq75W+3gGw4KrL6J1CKZlLMWCt+PHaCJljGt+wSVgzf6X2kMSeA
BIcTJ/qerLbJOWGfmxqbQ8oMI5O3hG/VOMHHc2cIWt6DI0zHJjQvVA8cQ/Ce3n5o
DGn0Lq0AbiMoH05/zmow4RS84AK7VtTv8GjUPPJu3dhqCYCLb0mSRDcDjxWhzi6S
LSFJxwPbLnkfrrsKwqEFEOPG/EVHpW9nu78ISx/tJ5HPqGDga/g8pBE/qaDKfeDT
4Y3BtrtbbrkA+QptyyV1oiO051JCty0wmEwOVC8+qumE1vfVE9Bp0QjO4ad9CeiU
dI5MZw4n0buhuNUxSLZhMgEgvGSyUJ/dtv2F2TlxgdMcxBOhTHNua3fsIF4YBQHa
o8I+VtCSZwQpYyCcj9zb5BlhhjQmHz8WbKi2G3CUCk32d1b8wjwWmnBgXdmmGPBy
9dHuUED6dWXRaxDf3GAOHrtu15Vg9zJkljC8WyW/E5xLOumKLj4htOhGR6yrxehZ
yabmUHK8hY6XEC4JTf9BycoiYfa6Rjds9pihrdZyD2eMdI+uYKB5XORsnjXAPtHK
zptjEpFt0lA8GZEWyDlCEDb7K85Cm1TLnVmRb+8L4pBe9CrLM3CETWfVvIA8GdzC
OFRFKIsGSsLo7kvR1Gy1zbGFjwya+S6I0TH8FtVgjEjK7kfDylqRjH/qkD05JRNu
emYYalkgKmFnXDe3WNAfGHmNJ3+233FqPUfB/RdxlougfJshjuSH1bHXefIbkmfi
BJGPylV2aX8OXkOEH+FwBjPciZmri8T4qEBlbKIw0oAm4GyYqTrOXANz6wYoSRHZ
b6EhJzo1WwbxEIUPNWVaw8RP2I0sEwuzAe1Oe+0xGoU223YwoXUquWz9f+RR627k
5N7sp5shNLSVhnsj1tK6b0ReJQ0ZCf/SGXcZ7W6DqOO4+PZxDbNwbo+EhxvyYoKx
Rqd8lrA6s8aL57sMEiD6ig==
`protect END_PROTECTED
