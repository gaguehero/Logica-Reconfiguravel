`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT2YG2wXNWKw4pPiwTaj5dnm96w2kXZY2ZOZhRy3YLp7egkGxgFGL8mMOcZQkEof
7w5hqDe8GdkF84T6E0Q2Js0q8Uava+G32m/kTZNLJPIv1XXjeYDKcNE1qv20F91X
PLJngt6ldvZjS6JW1pc8Y4eo5uF1iqs3JBrg2wEf7ubqEtOZbbDhIxgtqxv5vHGG
qQR3G4Uh6Os/ltHth7ZzHqW7JiltCS5YRHOiKeV5Za3ZBo/ZqrcXr2tr9ksTz8Nx
I9hjVzrQpVfG2saaOu05CnuS7fh7g34iY7N98iA/8igs42Ln8OBh7vcPacZIGC/z
fc7IRK9fs7esXBFhQAjmYjYSDimhs5dDKwNPonrXVjTbSEizazKEbb8fNNlpBgn4
2uFmufeS3BmfWfxJYbrrwvY3UXTzC7wrFIr6m2NoFfa5KABHM0IVder+B2+SC+Uz
ewICaeGqeyyJxCzoiQOU+Sno4D3wjidTMEWFKfPnM8Gx2xMZ50H3uvd77rPMWkXD
dilDMQmo52YdlpRx+w/EuL1ZBHkpx6CPQ6iQ2P4C5IOPr3MLWZFt65PZ2/1euHHi
056uNSUqiC/5Rd/fzm+bc8IjekJMmNZmK7M0c1RKbd0=
`protect END_PROTECTED
