`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+DrDVjE1y5On6NwISUR7Ga1a7u8Wp3IucnIZdCsF/X+Ig0gkI3Qg5ppj3cY8hB/h
UstHNEddDbSuiVrRN82nHrxqCOeVTLFn7tvtqHrvYHzLxo9n2Y1NqSoPC0OiHaZa
QHmj8KOCvw4N92C4T0x03+cx/dz/IM9anphprWRQFfRGfBNHUTqSiVrh8pldfcTV
WJwDTVFRRErOz5aTnIoMd0jpYh5ddNQjSriRnbMA+Scazoh9cfO1jTbcdB1+VCtO
XYDb/Ny101kJOCGyHe31QG29o4psNOlhmrAUwGWB0RjI/46MeCVjIrQn9M100KcH
S/ZEevq5o/p5EFQnHd49/ukxaXr+4QdUbOZO1Tcr4WyIsIXg7YHH7Br+vzQb5uqs
Q+sQM5GpmhEPa3J5Wak530MmW4C3ig5Qy8rcDPSXEcAR0wAau7ga+Q5LXgKZGyhk
CwJWdsJ0hZMVCP3oEqybvKrF/9mRe7R4z9BM+YLDE5Ch300O76mfZT0nAKWEmfKW
WLAjnS4hqiU2OGwlTy+g7x3Bteguaum6r+Ixgk+qdod5yjKwdtw+vg9Szdp6eVVs
h/rsZQ5TTUMSVer7xdcTJPL6h9/Px6zBcuEn0wG/40Y1iuaVdhj6Egps3tq1I+i4
JuWwNSnS7L/IjFT5edd4wOxrhmUEBGK9Ss3AF1BSbjjylMsYB/5PqYHkAT8r5x6F
XDEK2ha5jOvY0DAR859kPPwwKDWnn2JrFo5s55+WrPu3N2P4z37Dx0vrJxA2rKIG
fOJQMhzSHECY5YE6qwmKHJ9bcQHgNDHBAFz4q5D48wvFUpHNsdVD4uTi5lp0XCmY
HfvkBzCnnscBMJl8SWQSjvnGg5as9fRpi4Fx7YUhaFnVGP7cYvMoGdyYcDdZCtpv
BdeojWTYiQt8PK3Z5cljrnhTMLsxBN+KOHFVm3UqC9YTMMFwPDAwMF9rOM2tAtQY
qZTeNVQtCgvprtdwZmhAnVWRp6Vb1++ZEqVteA9TgkLtxsio7AgKdkMC3cweLg2M
nv/z6zxZg4D6rPutGxZ2dZDfGskkgOKkWLn1sp9utqqg3ewKGP69EWtpKCkGxfGq
4g9CYkus2zBt4k4uQgLqALcqe7b9EeTbRFoQ1k6OgIPCFlPfsCsa8t97h0rmYxOE
dFS0Cpxsa01+sQQ8GRMIhFoeRg0Bk2/uccavUphbXDfgFtLX2LFUeKemz//Hp2Dx
7BMHgmPtdjMNoU+bzQIXRA1J0gsL5FryzCfZQ+obtp3qh90spxkjDOFE91U/+DQ2
Hg+O2Zv2NuwGrTkrLrmKZYfm+/5vC2k1jhS87d/PVQdvIliWcP9d1iJOxvaM6UWT
aJ/ojBHUW3K5NENwebhd183k0L/4lvfkEy3LjMrpzHiABwV7reRe0a4A3A2boZIu
696ibjeL+2H7uozH86aiGU2ZKvT0CXEiPOoc9Y6KTC9cPysc7+rZFvemanexYIT+
hBaCtkME5aTqg3JiwpiY9HH1qIBPEIlNEXNn9tKG4PnFB95yMhpK07KxECAAUHlt
LPJbsBm/ZRWA/VaSp0HlK6jY7THiWiMwl9d+0PbE1/KhIiUj25JnglNH8ieG5Ku3
92fzUHd++B1i6p9w8BKrYO6WFPkxlStnGpUXViKWbGYgSVF22iTPz9nydimUczjU
P2e2hNAvyKyM6jRWqRazSzuuzq0hqHlQ2BE3ALlslVAwE92rZ0jeFsuGgaSvgXnv
Z4NvjnLNAzk1oO/0Nw5YDmKKy9nusFrDijbhNwsllu+4F2+X60rkb3049Gcj5bBo
anI1bicBE6G+cQJ+k3dN/LBWWGJdlMk9stTC+Nn78VyvOJw1SFPiiVnjTF4NmaBn
mZQyAcfuFUApuprT9A1zt6h5AfyFBuRIIv8qBBiY8yFVPbVHdNgR1CvMpq5UPgrl
VyZeTDrIDHIjR2d+2UPlNASjiDENgZEWuJrP4gBCMAIUyJ3RZWgdbveIWz3hzVZJ
Y5ttq+ZKVs4UAcei89+MZplmf7bHdOEmVTM2usMrzlmYbztkCzZrSi7UvSss2cvo
yW/y4WWx3AKr43iBEbh+fF/nH18G8etHBhCn5kDh5PPt+aX34CVXu6Y/DjHN3R7B
p9oy0naSd1LiPr5qDNtnbKs79a17eRIsJMPLhLhmie5ttOPIFJeg6lwMG0jqqaPp
kaznfghVAX8mM7v0PRG2zHINs4WClLJXDd75oYUd2cQFy0PY2FM6NmZRMyMbkPOw
5Nlp2xppOk6byAuc+Nv2KzBBUQUmxD7LtBPjhScvSfj3dAp29DeY8GnS3jAK/BnX
4Dahpod2WMK0fWsgUMzkLGKIZRKC7DTXV4gSfF4/Ld5HFueKEbzIdviAm+41kKYf
oHS+YGAWGEsYyFMKyR8v9wwOzHL7hgPG2r7FsI/2tNIk9rCF9fUZcDr5F9lSeA7+
K6F1SkDQHr58joQCsHeExLLWzeS7YRpykE0kh0NaGGkZFlnzsanTUjw/kF3Wrixg
T7gAG/pR2epKPK0hv13gP18gDS76INUHaEcFZrY97ePNV+t0J9jC1mL9RxXGPbUh
Z6aX+co0FX2Ezzb9Aj2PUmWSV2IpjlX7ikroy8vE4mQHBvC4BpDH+Ze64m8SBdaz
DT0jr3htmgJpuq2EboWG2mygEnUqqYxBJFASeKuE34U0JPqswOpmpiP13+lpRRcZ
rohmxDYR74DxGZ0l1f2Fes9dUjMxPYoFS9zWyfil16IVLw7+kt3+dRaAXbOacVUY
L/+upJsr2dE1WLG3jkiW20FtJj2UTjZDF52y2aP5zziyWlrDZJLT2evDDUORkQbl
5V65Fg7UVgWj4R9jSGNjUusBcNCYVMEBHs2aCgY5ql0lgckxdhqxiUWm7rQAFbm+
Mgycg5zE/M0f2dt9Vrg+uqJfKNIkpeW0s4kKvMdCgHzLRitFbi4VD9edtTi/I11B
O37UACbv0QN6dBGH1+DgaWyXPpUlLmQyqvEcrhd1V4G7zd6T1Ez9j72nshKjcer0
VUNEPfcfXX5x8BuiXu+WE++Nk/OgwCJBzRrFdj5hhAeB359Z9ssOQaMBTYiYWuPx
DTNg+ZwW57rCDEhMUavLZ1/OXGBqusmg/WRBAWgPM0cei8JXUNwhuCEA6ZGzDCqf
zwohPxgK0UQaP7fWx8BWM2k1ZxckUrYcFFHdKF2mbZewpr6TOS0fHz3XTjr6pKsJ
4wGysF+1EpaPmfCGDGuWRhjdpFUz4Cs7RZDoZXIpwuXF4fcD6ngdKprpxtKr+wsT
Pek/rkMTKzrYefvJK+RcWjkuCdwfv0tRf00IKDpVxj9q2kBgmGDbXE9ciYP8DXE/
OQQFO6T1gDcCCVO4WQezm7BmxOmXdGzmMCYHxuJpgkyux/NQjSaSkZ/VQEF0eUUY
tS7QwCKkGxwjfFgZvwGKuU2DC/oJHiEVWEmksb22kldSIE7YXhqhl0gWD4K0vK4u
KTMVN8eGgmwrY2e+CqBcnLJO78blpn4M8U7YNQfA3gAAP90qklNqswif5w79P92h
FZ8/5RRS7wRUDMRSXL2LTRBF3ZOSlrKeZtn0/nobANCrXpnGYMYNbwj9WLH0DCzo
fBhKJP4unuCAqbJjdFgtQE+tw/JLoTCH0CAujTcFJ06P21CPhrir3K6UTfdGkzqn
iSyDaK1pZQeaq4vrXjMZr9UMt5J0bhNwniwx3jstKKqC24KVSeBuyLG/LplaKey6
ufFchwp3rIq6M3W+SP0SrpsW58AJU90OE3GtTq03r/0y0/lRpjXMSctlOS00saJ4
f347vp9rjDSNX3PDrx2TdDwHD+f3xHFXo5418cqAdKJdz+UtXjcGDLo12F1aQc3P
6YzsmgxQ+8DFRrZ8Yu5adf35ehMAcsGmFToCxNyPA1esmcKrL4760a+9P11E+U00
XrifCPToQn7XT/XJ7aC3BXbBauJm1m3nLsFZJ1HtnSmSyn0AT4UlDQrUVo6HD4qR
rETv7UFx1iflUyae6xIPJlinZ6R6MSerqh3UMFx/Orlb5K5PSXG3TmTjnGq/kSCq
taIMkhg3S/np8252bd3AOJujBwmcF3oUr2zgQeQIMe8KJoB3jzPm+CWU8DuRxxqq
1qz+FXFRpsbhFpP/FfHgaGcXuf960QPKK9aNQPq+UAHiefVC+4aTGBfd4EbQUWBy
JtD/ev5GT58D+nBO+GyUfa+2qnbWjL5nZMaTHFrg1vhOB7eEYpnMNoikVfYYQ9iR
lOO6SSCqKpgUIHZLU24LpSVjaDvLlhWJRvQU4TGj2BgdAWouox2CB4gMdvBGZO6+
IOyCqJsSevevhQ5UmAlKpRFlbHY5H3ddKnPdgFff0+QwQt8VCzYcCydrVP9unXye
zZ5Y/mq+2OYk5RgERFSS/mmcaDpNJntxf9KBOxHkL96eUYCdl4GdmV2+gwmN1IEo
QrEGrDXCNeiDsvY9JtFvRDK1hOq3HgyWzOhXYN1iWLgM9ZfFaVRqM2/eaacMR63n
pZefOuDe2UzrgCu6qSZzBn1J/XNr2EbUVKWXc9oDbXLm0ARG5hDcm6WF469H2AmC
JTr/kmadgrLj9LS/4gNpvJNp6R6Fodg12GVsWx7QC54FIBynVG7+1g5eeU0AynSf
g+sReafC3+XBalVAti79v+Nufaq6CYu77lVCWvbB5hs9QSojYmzzyueK4siqTMnO
05xQN7XLKP7Ik7c5VXpIJscBmN/83QsUlBkjLzEprhmfHJ+F/ut3+u07te45PSmZ
N4Kqbcdw9mW722JE2iLx8Wff57PIk+f/J17QiH1IVpIRoPQyxIUuEepW/OKBhtyY
uAWm46o5ZSKjIf21YFlP3isFam9oC+lXb7taBKyuzAkIfQZaQpl+szvCwwnmqzuI
Sf6eki8DWtlfUqb5y0SM4PVGudA3y3tW5mWIAQtjQQz/J1Uh9wIc/3r41asXw78d
d3uigyiylvluF4/KY2FmDszUoOpqAwDabfAkkmVOfUKkUjiFni/UyExTc8J4Jf3t
oduQPssKXdX++in/cTEuN16x/9rFGj6SlW91yxHTXN1oq8O2A0RiSJnGI3DjKPSz
oGR6NupsJCQ+DiGYBeeDP9ZeUrqwxfYBx5xcLm3efO6KQfRp7Gcg3JqVs7V2GMTK
WONtShjYdcFNZIv8rRX7V0EHiZa4nQHXwAfK19L71MLRem/pNpuInMqnGqfBSAvY
uL7+bB4pT+yT/7qNuJiS+0ibcRyUXzrREwR0Yjj09ApwMh6jFVvHSE6xG3mUfho3
aZj5YNTLD2Nqm4NkQSgUs+gWQ+dLQLTWn6Jt8T+7jeAqJQ490CnewaczeXRsekNL
zTyY2jg5K3zSl2wLS9a5/BEWdo+uLyBAK5zETN+7ZAxiE4deZgmIwzYa6hVJezDc
deZLSiorz6TPBhEj1qX8i42/bmfvaIeuRA/p8C1MHcAx6PCJC8gmQxYiGs27u67u
RTuIhvRCzpQj1wSgMDTJTcuzVSR86eKxiC4wtCHqUQigix8aHjgXGFuLnEAPDW5t
GjwAe3aGc4XYMMrfX/dT5OMeLvhkFVt0W6i/RH3jUo+atfjIEd5aJMg5OqgD3MpR
D7Ef1eUKBrDJqFet43bTiMpAnt4p9GT5zQFovlmVU4OjxdBWc3OBkEXdWYP5cIYl
ilGst72LGvUZgIwk0uSZTQIWks65h4aYyOoku+lbmu4ugIfbHeJET106uoyFHz1u
lgr0VADQcYB/HAfgICTWZFrXp9Y+1xdMAWY3PB0qrJ0P1RJitlf77vzfF5J0N6uu
YDa5XbKyMOaeDYKDCh+1scAdZvLCReDzVx4cJqoJI9UYdFStzy6v4fI+N4FN2ig2
1KpY1rIYuef2RTaQ16ASJQgbg39ZsUOuUq5Lm2blCUfpc+VnWo8EW7N5+DOjqHsX
n8vsmVwmC3+Ct+6FUj0nipKtZIOB3vF5QFoB47TauOyOtWe1/VVY56OSrODiDUyP
rVlOzND8KnV2/Et7lpC8YYIDeHLYYoot8MhpbisHZdk4C9WgHAVnfY8Dp35L23IR
JC7y0Y0w97gffpZ88kTtUll/2V8EbTbbB5C3U0N5XoN20ltcal7sgkZi+XZjhpVr
AWDaCD3g1Hw878qpp7GJbzfD4oUHwJMedtJOT8cos/OGzhzY/Lp3uW4Lp6ezJh0W
JPQq52PjBLGFoYpbL+OJrwEQfHicsPtg110m4uy74kY1ZuIYwjFMCOk8No2yWfwf
sBYMUdlMr8XlUqOuZOfbITyf2Lici5ZUvLvnnddxRbHwVWvEd6vwThjnzF/5JLeu
xMex1YaxJIoGHKYXPJqaNlUJB4reCiGUbzFV4n8s0/bwB98imd2VRajmwJqu/xBd
xOynEiO52Q7zgI+8azCvWgjH/RObKPzEFQ4YlLowbHgcJhpt0K8uxgGaDjX2ZtXY
mFWZzPIxoyv6bd1JdH4o1dO5khuVUu5D+UZjn1TIpxbtMFp5pdaMT7UKwYXOLHj9
/1WQx2kO7ua3e9v45qWTMw3vLs5u2k4LKyrObfXUVNimegsG45WHfPDm+Q1+MhSR
5cbJ2xoSpwwpPWSqeYD9t4skE5+zxjJoCCjrOQffTEa9iN6tOy2jQK0p3HaHRFxO
7nwEWh7ssvzb3opKmeMWGUcJWJ04Ek2B+tTKsQgYLMrkzRJgF+DpFhSVq5dFBIB6
uON1wiIUzy0CE46jGKB+e+bPqD5JrtlDBC8m1xbEYW519IGtroOP6Lt4q3/ckRDx
JMvEFlUp+wlcUHcXQGwdi0zqOEHufvOStHHOjqUQysrzcBbo4/MQiYA0h5loLW0T
NbNaccXjfvyxPZzYCiDfEIBorrYVnXJe3/dEBpink2zqok4faPqUyqdv9bjs4kJZ
1xbckMYdHf5npSUVtiG6xZq3yawcOVpn1nXutzKl02gXWQWILAxxD8u0moU655EH
sHQUp6nJk9/s7XI+UF6GaezTkZ7IBm3fet2rNpKIinTDWpjxmS0br8dI7qOksn+m
UjANG0Gx8GwJxN2T8GZBWI/k83Z3tQDSsXr+j8BWOwqowTWpLiaZqdMWzpdqp7tW
7lqLhq11hHPd6ROUMPST6tO3fMfA3q0+zf88YBAOVS5g7PPDsBcTZdlqH14wPc0o
jBsiXCnJBqQPlNqSaZUFX1EzkQijRdbpAcAyfxCxka6D7vE9uqFgz7eTsGaiiuW0
KkvBJi9eoA4b4yFgm6XkOl0cBsrpsYGD3qetnK7VgMXr8kVfRKdADHi53RhJdviF
nK9Bh1stw8P7qJwq9ELNiS90dOjV0dtawzubw65J/bpSKlLL4K6TolzF2x7TZ1Eq
LgtIXshrFCg9KO5OHtUFFvL2FLnGre4XEWiWMDs/qz9lUT+jJaWouYw9VziQoQ3W
XoBWKADa/1Qk10B6VGbgw3WMhXotrLjmePhrJkO9BSqabgdPYPWWvd9Rlic3cjiq
gtj8LsMMpTnj7MKHF4g/wzv9gj0YLFrSF0C+x4Ir9/5HgNjgLwrn0LcmjocsO5KM
gXoqMorXOOvEMaPntRXInIFZMZ1bduzh5Le68dDqlCTKYbsjyxPGn2Cjosk1DXmy
Vkn2TnOjAWZH5odxUM4KAdtyEcJWGJHZethoWt3iKjA3ywH9TXSHq7os4quwcw3B
Tq7KqyL57xqWwUdqgDWc3EDUmsVWMqEqVY4FTgeVbGfBgyn1kwhNXmuoaGT9uvyK
`protect END_PROTECTED
