`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7Tmc5Bfp+c1LED+hXR7yX7+Bn0YfhXJFme/z2Xo0thTzE9AsFdmcz71cyyPWJ9z
ewVE2IiG2C/4MXz+BOCIf01+NC4CTJyoQ1LfIHoVnDVehyReOgcrmRcG9NF+GT/1
h6EtokbgxJOW1s5dKFSzFou2OTxGHPVUTkIWWCfjaKrW9N8DQZEKIyoX1sZHDCWO
a7IqxCaEs1LpmqYasfu/HT6fp4qOguMYw3jQn4YAL8x44iG0+rz3ljKIA0NiXG6R
NCPnPD/FAXM7JeFocaVu+CzI1G8HeSKIkJkFhA6YhxZEf3hHiC3DRcYSVnFRpwgO
J3HRI8I5vWadxEKjevWWgLzZUdtGgw8axuDB9vW+O9pu2dmxxeLHeKGtUMMYFn2d
sac9RU7vnoLhzGHYSzVhN9dKHzTy4cw3t/G5tv0mE7tvwu+zR/7ORQGr8LhFWxmI
NeZDy3AtMWTAu2nb8OvK5f8M+Cc7+1frmGlLxyS0PRlJjD/ZOPI9sI2iV4X/W+4z
XTcAu16J+3FjJcoeNqcw/a3AzXdKPjUW/3OnicGExlUXcOgaejJ/lRjJ5xL8+Oyf
VRS229MtYk45LQflTHVQwmND+GvGHpfgL0HeAKSQQ+7BlVGCIaTzjL0WmBrY9zMO
8V0F3fEW1NH9MitGLLKnaDJ/Zs4Ohz5tZyzCT7hC3VolbQT/OdJpqft6O02q2V5f
U8p7hGgGWJiQYD5JN+8XrhnQYpo/ViCcTOWylYW1orQ=
`protect END_PROTECTED
