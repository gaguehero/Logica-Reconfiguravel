`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o9SUWcQxvE9V6f97AmE1epPKE8hptgLjoNgfVJPyyS06fLKVv8vKss7uI32JBDfT
9tQSIjUrSzgXWPVolIeyNQjKTgpmAfz9aITna5vHkRSQeV9jm29pCQHVd1mRTrrs
qX/whOslJcHci5DEWh3izsChZdx6uy5jxHcAZn4PUMvdVj3s4z9pbEz/qjuQPdGT
nHb76OGjTTiZM/s4fsPDfzAkbSoLQKqISuvR39hvXU/acGZ7f1sZxgpHiwUkONl1
LOneHNZX3XwNf786lQGOX2MvHwUaHEFw3qPB+P8IW7edM62VSO3WNwlJ2mHdUfRX
yIekNLZU6ABlLX1Bveir1BmIBEZ8xBpN4bWAOCY6D37AGZARHZJ/Q7YRCK0Mpt6V
oBu+V92fpeJRQbjAnFrs0mzpoTG9kE1JUpsKg6pO7nU48MDzf+vWXKJzqY81/4CC
aBROxuVQWX6DGq2RqiqDcyJVIIJNsSut8qMVAlqzxb9PNC6WrskrNFxXpUKxhkfG
prVasu7F98ZRb5kcBnrGsJaae9T4CH7iAwcqz+3busxtE1iJctkGbgl7CdRV9CmP
jm5tAXFKKp1ljByZ2TFlyzqFVbh3w2fiYoAiYXGYwE8fCSCZo2KYtALLIJyXpZEy
D9jRawQDYHbAIzZiRagKLahLllb70GUCriqLG5Uu25U7dVJSSXcjAphKZNUgyDnD
LQHcco0bsMYoO1PywqCozyWg8we9wKTSI/1dDnLPOww=
`protect END_PROTECTED
