`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvl0GVy0r4lr/Yo0DzRNWpDMcktaSaUrJg8rWjfi26EV+DRpr+OuadXe57qkTFgh
6QpLHEqzQBX97cevxbLWAfToCr9Fd3drNkGl4mI3hP1vFqlXmTDYHkrhBf1FR7Gw
vUxHhaU+a6k+4UHhi5JPkoObInNVNyYKL2T6jl8L8g6XJ1OmkT/DtiMoo29h0ELX
AUcSOyGQTencxF5z7RZensX6xgMel6UbMbH1s7o22rS5scHQukLQ8HVI82fClaC8
hQw7IIHbo+4HrGpylerUDc5bLTFiuqv8B1b8IsT2OGlZr3PtwW4kpZjgJBgKsz9g
/LW1AisIugH8GsL5x/+58DPsUwnAktsmFUtZN0eTSxdlWVI81/OWGI/y0bvqI9kG
BRRfWRJxRnertLnfVJI9nT73jgYvichvBsSpwqvrEeVvZFOppqW+vwrTqWsbnOPm
+BmrpC+pIHr9DOQl77mf/t0ZfeDtTTAGjxJQyVEs4YP2sqZLBxgLHHOiESLp5BXF
pyjA+dNvkRzrHW44iqD/Tk04zVRYwkcGdjxSbQXkQUX4gXvswIO0eLiqW7PaUS+B
98DQ+x4/utBw66kwm5BDwSHtmjG21+4SYQjzZztwvv/73rMH6rd+vg0MWr7LhlaW
idcHqpTf6ZeApCTeJdUJ7eA+KAJbFcVgFVIZcUP38BKHMexJobMN8CNI8ZiyUw7n
`protect END_PROTECTED
