`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lfd4DcvjAtmd2cAvXUbxMOCU1vM88TJ8n3EJ8J9X1ySLyrjx36rHSNM7BImS/4l/
PTDcgM/Z8vT7AS7zW+/tj766to2TLNVLlUvkVa82IO5g+umTw7qJ6MKvYpmafbCE
1dfnlBWS2yH/sBsfizCSDruQL3DahIAMPU7BgRvGH8+N1pCSXLshA/Wh93xgc4z4
VW6u3MoLBtwjymXn3ERJTIlIcg+6nHkudTkdVV/LH25vJWCwPRqAHEAlN+3HTLim
PwN5sWQXtQ2VpLxws4TDm5xamFOhOSbqeqaZdF88WWfrpDNaOOPCcx02pVL9D86n
Z8lqkbOkw/VTZ7cQHEeMQowoRaIby9O/syUErHHhq5oY0ZqwdDQwJnazXXCrujWX
7YETaKVg9ZSdG/a/y9QQ87ZYz0LFlEAhkKCrcXvYjjONR88uHy2O37LjF0ICgEBC
9ZJewgv9NfrHh2j8ypjmfTskTvfOTB1m2Evf3WmDKMpe4W6VV16NP9i5KZXtUky/
qs2Xpk3/pnNVlK+W30f8+ucjz+R/zQDaF25JwW1R0t3XKJwmqY9JqoT0nYGgqRvU
GCD9Okn8L0Ys3jGCvLsfhKMRDnRPkq2cPcW2eFMTCrrYju7A/Q3al2OSVoh9CdbA
pIAtR0jsMBkLWaNKIGmNW9BnBzlJueZCSE6WjfG44bVEivrD4Xm6TND8x9igC31u
GWmRxUA0Ddkxc+aQ2iqjDcQkALsNOZvZYiYL4hkir6Cf8A19bUi4CoeDr9eklySX
4ArYDjvkBQtkboO7qHFy8Rt4xSn+HlK/o+fbMAB12Pc1cMQJTyUiUvrIq1zKsdAN
Z8WzJOAgtVzNHsa0tnOxG/BcuSwlG3FyHWImbX+1+Xbnj63rh1gk4wdikn9qsBgm
7U0x+/OGw61xyVuP91+LOKEjujgUcuPOnR5THDkyX0IA8FzY/hK1qz/O9zElyI+G
62qtSBXKV9JzzGU0TpNabaAkjuQpS6rfvj1Bb+RK2mVGDShJQ8a5HUwLYwsPLxOs
Gr2ao3/nI8whOSDdPicpMn4veFkRV+oN3HENp2tG1ei1sMTNMZaRTUrD6d4uOonZ
hmD2X+0UQvNXzCg+S+nlWQTQekxXQRMyRf+7sStmy8WQV5THCPJn9i7uK8I0Shz4
Xl0kbPkXuOunGFNA4k2jmewoUumq9PGkSAH4FhOAnHAe8VoqklfpcPe5OmNdI6cu
N+RIplnazZP1quUQscq1oWvTeJIsVNGU0b2oG/+Ed73ULB8VKj9fh+ERTumXbNdc
O0P/dEm/DOZi57yEh3wHB2umGoKm8HsjyJr6WQ6f1VGsOOJBFqXG4lqawhpz1gCn
SyJruqziEschWNY+LAOC4RFrNr3Cs3ajmjgu203z057IzDJS07SGY+yDY42s31np
GfNqol3YmZLQbkgMc4LB0XKW/05LCLFq55NHMP/bgKEr+Nictt/MYxshw1waRRro
XdsH72QTp0gHUJgbKPl2zv4khDPPyLBu5t8MztyCs65K40yWzzbyowV/NdC5yFC8
XRyzbf5o2gsRAWW5ufCEJ3gj7WdKlZPkzsfy+Q2du7LuHitSOiUP7/U0R+JuDUt4
KTS+DWWqYk+0nqtYFXHfltmclJz3fGAV9G/Ly5qSDspLPfLBXgzIs7+Dw0IWZCua
f0igyTLp4VnCX4Z/Pgv5/xzJ0C+aXCb+3BuviheOBKUbQNmFi63UNbHZpTUQ7/V/
kXb+AkITIlpzvp65lvb7XlKMJ+sxqu/0nAlKy8x1SbapcYeq27dsa3VZwHjwPRsm
3owvN9c/+PZ9kofVBYPOkMxmwNoSUXRvpX3lSc0QvMjIt+nB0TEmIuadnVS9KDt6
GMtO9wNL1WGA5JgnyQ9IUbRMb/w8iOmuX/LNU3iLyRcDiCDcChS1g/ZjElCe8EX8
1yo3JaEA3+LypjgwewD+Hq9QxfgoJ5q3Ir/n/4mFhMyg1SQS8lsf1r1f2aClkNaf
77yx2RQkkf+onevLJLXRF2wn1D9hXk6L+FWrWHaA8oaB00z8NhxCo6DkSy0ggdDB
`protect END_PROTECTED
