`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHzN0TSOhm0Y4AyKd8BpV/3R/2wrvEcRL/Nie3FMdELXqBehGH60+hvfcCTNoDly
yAwfZYrQOdJTZ0bPvaTDL1YO3ymxDgmIcdlRDDLTlI2WiBkkECSDGiCPBo8xIlYC
6Nd9QcYC0gQCOHHvQgt1pp0IW9XxUxi9KrO1VUC8UAhnIZvvCYlhdPHSFlADQEIM
juYLuLmsLoh3vkBd96+Egbr7+s2JtQPeLsXvM2XurKeTyqRnTEFmT4XKpKbo0O67
6bkvg9TYkO35mNG7RZIazrlFzYw9S8bgo2wK9ED7m8UGTs38IjrlMFZfCPvcs4aC
hThH0pScH9MmqolIDr4NIUWgY0rbB23joZRLmplZoFmxPvyf6RgiXGIn+6ThuT/3
+0e4Gz9FGNMyh1K/RGOuWmJ+PeOUTy/CDyggxDz0JZ/n9b28tCHPLyA0jxpBBYEh
q3j6gMlXuNlwXHKO/iJIwHnFajQ8wEkw31iImgA37c123+p8faAkU/zVd8FOmVAu
czmQR0x0bECqxi+AvOsyGdP517hM+QoygMtw7AuwiF15OkkOVIU4mYbxjSqyZite
Ucu/T+vC0/3A9amJx47vjTEHSrVpaGoGYXuGrcPKqF0=
`protect END_PROTECTED
