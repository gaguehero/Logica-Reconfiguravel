`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTr/0QbLJk7la/IoQwk1qnuZdkFICXSms+7EKfMn3pXUT5ObQRDObjRW3A2p3RHP
DzHJnk3Pv3FQFHMI17pUUjopoeBri+wpl84SwRyVWlT7Xjrzb/4TJe4IhBUCFmy/
7pQ+fdLDdKPOXB/V2zzzUvB/0jSIcV+x7tjWJQSA21TKazkiEiF5HnTvtMtG0V34
LtVeJbUoYZdBdm27NHVzxuOaQJMjJ5JyG5DSt1QrY6Ie7HBc9RW/K86iUnnTxEFo
Xz77/TLUfjcRBsRVyOFazktDsW5e5eXOmHW4cNR6DtsA7MxezhiR7PZ+qunTObvH
VwLGJYOvZ2z1TQ7dGqDpyG7WLIIOB/3ebrCyOlBOIHW570+IQXOF4/BuJpNRgewi
WJlrvfpmp2l0wbQn2S+gsJcPsOMqVBFo26kA+jyp7uotYw56FH/1aLuexAMPACTp
4H/2pG9sX6233W9/u0ntRaqO3mDHgg6mmJ/G6+vKSYM1lVLxdw6eodHPkB2T8ZVL
hR4W7ggoJm599A6ebYCN/RlqvgKCz3c31n56Y3yxLnjJUVyOMmvLr4XkOZkgZ4TR
HUZ2Rw5cZjiLLHRB3DtdbOrQ449o1UVxHb9HgimETjA3NjAwTKhKMOeeuJ8TmyAX
dukioMo6hT6/K+5St4xOC05JgsovmCUP4kr90BUVGvjq0Uu3wJkp/pnNJzfaUiCD
u7z197UI4uiuDS8UjRbxjhFOWMuTVJde3gIUX+oFQHk70xzjiO9s7AMtomgv8TXD
NH4RTv299+oQec1E/ZrC0kXSoKsB8r43ZFQcdxpRT9Q3H91ukr/JnMkxnTDTyx7w
TEC4TR6x8ON96pLoIfvTjX8OgURh70Hbe1UvwANshyfAcgvbNxmP/tBh2yzRQ+HZ
uDz8pq8kTv/Y/6Zlh0CJIjdv2tz7ZkKIA+WwoaMQv3r9rnOyC3wYJoEd5fIyOdv0
rg2yAHQXmp3MlHEpGCR3nZrU9CjOhTqqdGJWFDqcZucEprqPa6O50+JPF7Ozc4kY
efFmQQkqThRcmFUTQtnH6obdKKjzG8VsjSZHQ9f7EvzDDUn+mG8sx2a2gHtWBzbo
WzSH+Qm7l5YpHc34DwfTR0LldtvzjL/zB4MmTgwcepGFq2L3NJ7B4ndBdl4DAcFw
TXUFXpyZ/bKBlr5ioGX+xc6bcy8BIoVwsffLZESfg54ymfWdFTxMsVxmY1UxJGc3
QarO/oA0B1+T8ScoreKdRNmZeNBwBsYJ01l01kWBThSCSrRaArBH9y3mKPt3cESL
6zsEwRwTZhDo3N1JUhKI+/U2Rp6Dg6/QR/6kGxKB2K22enHIMNqoFElD/omnoKQd
BnlXZQveMP+TZMkmVIGDsNCv9WmQz/qp7jwz7hPcegmQxvSpTa6/vOk2KsVatlmf
gltzfd93KNcmvu1mJn5Oe0mrgaVO5HrivhSNdnaJVWRl121SxXJFwff9kmdYhG2G
t3amGZsKL12UAwYgE3m6OpOKdAfwUGyZhgIEra8ullmlLDT8jBDReqAKK7QbXvnQ
ZCl4aJy1s2bsrpgeIJaX28W6+AzxTkTgSerTiggxyWczOpoZ+ETDUlkG5lpeN3RW
up/TuNqS3xQ9kr8bEe+SMMojshgAbMCYMPXqz3n54KhGpEaKGsL3n5PIYYVN2pRN
/rsmFFmEKPG90ggexvKhmVylG0pfTNpUwljYZ637GPK0qJGch3xtmqLWToVyU3jq
I8nsMdP/s+kTZLyG4m7EC6tVibXVYmidrpUTCfeGCjGpvaRvoE1J2FIqB5zhZwzA
UDqiUrMgN6JZ9QYP+XQA8EzbO7rZ/rWgiYrDcrdhybUuQpGs57LR7oksH3PBlnbs
oiyv75pQ2cDW/HybN8LVL+mHy5jYiCI6qK5siH6zC+5EMtdPjBU42DCEcapW0ULY
r71HUcVV/jK1WCFi0o9ZGm9z3UI1RFFA5A6LaTmR+r1fs/WCtbgwd2nNyMT8YFx7
Jo1buUavErlxokOdGtf0KXrbKpotagXU3BC5VusTrpP0OWIrP8z+HHfh9T0czf1T
B66ttLwhlM1q1nGMI+T2f9lQlcmkNdLIPaDcb1+G4qFxtPuh6I5Msoo73v3znM9z
cyQdAfNdCPPM+8QeGLelXuuONDnvnE/mSOnjIMT3DLWTLUOm/jwLASe67uPXGxkd
zX2L6Cfcu45N4jevHYasuqaocUD16rIEurLANwJUUjmHOOc5c9xL4YYyGzAKRuYL
W6ljy1dW/vUBHkU1qURl/yukvjvSu0unWjo/lCih2SsndkZ3UiAKCByFSpg+Yg6s
uxn8KrqOimvo7fDG9wG3neaT15yoXAhENLNrb3LY+H5TPs9b/ZHQvpZCL56TxOGi
YBxG/ywUI3eVhYXgTL+f5uRB8VzcX23OkxGsl0PJauvTMx9zMZ0Fzlte/FeLkZcl
m1rc+jzKAMyt89DSB/4zOx73PSxgqiAhLJoBG67wRbE5e99Id0RciBvhy4vjjvb3
ZrmoU5U/srf8zEw/IE5am36N1c9CPdVBNT3Y5UIPzWW54kmoWXB7abqbspDXKpWe
NcuY0dO+BmzMMENL/iU1OD3Mwtw/KMv3Y9QezA4vcmEc7wHaiBXNczbRDOzNLUbD
OmtV94ic5s4NzTHcNhaiS7IlyCOaCKHdZRXpkXngNhl3zgw3cOR6ltk++eIesgEL
UHTOHOW8DpV2Qyk+X66D0JMukLWJJK+WQ+xzoAeAGgNIfv8HPWegwbWsqC9N6y+i
KSLBRr8zJoRI1xHK1+QiiIsUrXQCK0DUWWJ6/NYPqZ4CLZ4xlF9onzUJ2rfYRv2Y
wh5hM3iWdaTf+8Byu4/vm6gpCNFwbIGi6EC9AS/g30md0XxcfpGOh7ljH/O3X19v
4d/Daa6SA0eloae+j2EFxHGtpC40m/oanC8ukm4Oq/vJ+lpf3OUMTiRZf3qHhspU
LHUPe6xvQppCiXvEKcG5DkNFA3VCfGxgezvN/c2T5zYUkGqxNaHA9g6ai4E5p9Ik
QY4R9bWvkREJ4BeeYapBC04vF8MgUls0SsG5JyRTqeTqSe9ugZebO4+RCSmr4OL0
1N3beX+QtW8gbLRK3rvFV2vCrhkiVhbRPRQdzAjbkiWujLFSu/c0HFz94B0i8GVd
xEfXJ6gLRSpKb8NmohwzdK6L6NEqwaALL2sHBh5IB2B8Y7T0F8faEeCSL/AufkaB
E7mbVp7uS3kmGfBzlihkyKyyr2sZBu/AFCpNDEOfHOgxPEuZUn/15laTqCHKonw+
yk8HMsfOq9zbq/FvEg/DQ81QeJcuDfZoiEDYCX5kTIHLKDNk34/ys0cKn8fM14fD
0GR8YtnqEacT2YFe1PN+Q1yDTW879IzJdNciY7TgItsryrgEoFjuPPp0IzG4eqKS
usW/sw+BMZdhiLNn6tqJ3gkgycvH17R8hzvUlRlDm/s6oRaNbO+cAQyh+8xwGrPz
Arg1gefbuZD9kINVKqWuvUfLrII5Nm9vJpKlezdA21R8zA8txLSFYC7iHQEylnXS
v5BMNv/7m2fSQVNmeiMZex3uUkSyTU0s0eTNl6zqQ+g0olte9QZwP7E/PF5fNE/f
IBQwxZ1qv2NcAGHvORFM7sBdYI7czPVgGrYNjNf4N43UqCIOCorr9u8JIXlAT5WA
8dyIrs3QAabCOr3Be5/KBr9pOw5d9tGCKHlkj4EMpHaTulLHHNv5L5wtC3cq/Pb5
SbafQZmNE8CGHSWYEH1UnqVAbVSUqnO0X6sRjIYLszFP5K3MlBLOWkttyHsI8Lys
6Jr9y5ybo6xNqCML6k72YgbW9RO55dUgKTUYq4ko9RzDUssghFGN3EjEvnZt3Qnl
wHzMwC+Px2TnBAo34D9Wx7xPomVu3U2sCs5ntwVt6J3zEavQOSYL3BZdgCcjBtK4
+dxvK6n+YE9uZduG1l5QkbKoJjFrEbR4TjQXwEi2j3pC4aR/dZ6i9Nmg9Tm3AmF+
yHkg/Y+LLrl4KRM6K54WqS4/YB7OihwRP0K46fGOgnQ42iRKhg2X1LGi1XflFQ8E
OekIMRIWhZaJDjU0G3aNmOdvFnTVHM1N8TlmyK+/tql/VMHj2tQMy5ogJM8POL4W
MBaLUyECWqmvCqWXN9NYtULlBuX795WYYCyyyhqumbgbd2CX3F0lw43qoOdEwvWI
RJMvn/DILed8rd+6/SqJ4Jebap/CIEMSszTrda8cX2e7hMZP4S9n/7J2rZok0nwR
OC4bMayigWyFQf7pJ6PRaowV3+/iIGGYx1OhQVw5aea3Tf/t1AUnwLYdqhOlK1lZ
hn3BYW34j7eEWvzSS0sZXkEodwNbtLIeuV6zdyD6aj629OdYGVJ3A+04Z2/HZROR
hNP+XFtmbZ08YuRUidcGWrM5roxwydk5LMOuJ5oAYHz0WkjIDDWn7rz/4mshNKeK
WrSxZhwHkmIOaB+cDwyNqB+AycxE7cTsJU9+axcq9BC2dPFik/qWwl0RVVG9hjTJ
oF5hGsc3tBKAGSx0oz2B03EjJpbIRbPrxVGDoCaS97oCHqcBUJ+EpYh+r6KIRay+
IJ5vVdDGCRdonshEg2kZFhXr7z4x53aFHvvFvAYN6T/77MxPkR90TUCEtGehP3BA
tkU+lntykd5RfWLqNib2yDepECaYKaHkEdx9pzJk0a2DAjO/Ds8D4rS1PSkucdpp
ZMNHS4tGivSX/9eQ1qWrSpr3MxEfFsEIbA/orCU7IVLaldCv4eK7hlo+mjHr74k3
XH0/gTtZIX/bNi4TanZx4LhbT3Ro+BnJSUNPL7CzAR8khkogBqm211DVs9/E0aCe
EoqdXMSjkAeDHB7tm9+2S4MuijfbidaiwCCY+7AXm4/IxwCo6UxmEhI0etM3j31I
fZnyBpjTJmYqZydYcCtAW1WrBQFM/ARGPRkGDUDNaNCr5U7oEe6GSM9IGjsxdBqF
Pjyvj9wkPe2d5cjFLumlSWdQfcNwxFRocH/e+cgTvkx12e599zfiFDsOxCZrGfzn
JMsS6qgz0SOsiF3HEwh2U++8UNILmWI/YdonHaWDB4Pj24d/4CudlkkzKhz4Dgh5
c5kYmmT+ZYYCb14zcHN93Oo0eOCR7BABv69qJ33gEuXHICldNxyiyGg7Mcgk6hsy
xbC+U2wP2yJRzhBDWiK5IkE9SGfaDysYFtQY6UYaNKgS6lN+KnMLcag6PgKkikAK
T0BKiX5iIsgrxuHSfRpBqDtbsnYigmhFXDJVmvRuCLoVoME/1FwzMNTexbrTKwf2
iIgFRtgcKW3wwbN2VPbcn6esVBMV/h5xrbm1KYLoFjCRY96Oag7O2OQTjaVbRIhi
xW7mTzH7Sj5/XvVM+TEjlBZQWwNsawF6nJ+gjqg48282sqKEVMPIWSmNpU6t/lO+
JvOXEsApd/j0Os+ZAJCf/KOc/tIHOXiUds2S5MhqLEWgu3+W4a+EAwTmm3zTCmjK
fza3PAZmdtg1dBfwMstDj0CBVOyxwhwDuuO/xAQdHv25H0FB0rgHSiU2GbeN5AeN
soV/2PYZo4ljrQBG8NB7P1LgpEcOQY1TUWxLAFemF8gGbkkhstHW0ZppWq+z32bh
1JaOPtcw5tNBlLXzkLQ1+WTAt1/LtMSa7b48rXN4BJELw4oesETdgSzrSoIxUwVZ
IAk1DUH0Gz0QCS2GOq1RH/twUNErOuApeOj0Cbp1q4B8Rh2AhWxk3nTTupc2YyRF
CYILYt0pmjlLVxXOtIenl8xVC6cXYqeQ8TzcRsERXj9wBa5ovZjbmeUEAPh0G1RT
BjvNpNrZVWNOSpP6A2llJQvpanCZO/OCEjCB2rI5xNER/v7tCFrZiZOt4Kxkm390
PmkOupbCt9wiM4tWk0UQYQdipCVLjaEuTJufB1WWroRwOFQ4DCK94OGFIye4gBsC
1KZ56fLS3mVeXVP97dxvxIHp9YjFo0LJtTgxgxWHDnGAhl6Kuxmiim7jhXq2xMVa
VO3AfPqjVGlV1p4rU4qMYPOb40021aOt5uPrJ8y6Cr2p27ECExE9BBDyN/i/xem+
f8A9rllfK7QOby3gzB26A9dWhRxwy5mPOwvWUF3hvLaoPzhdr02Eq8+dwUBtnOiF
VXTvb3GYCxlvdtFFV0KlN7DogymjSZ99hTFWcQexNvoXyA75zdyfPLlp2YgVpfsd
vuZFabVvb5AEAz5vbEuM8VwVJT4vCGQg6dOSsFy+EdW1ge5LTJcoSsb21Dj15eOR
xIIFgB/zLL9HSMxNsFg33RCUcIAENbhTzYYkBKuJVY08NGxiyLXwUy0oZ7fWFw5/
ioOGlKFX9GZYYyhNhCeFljUo44vCRN2+7erAVWpeEU86AbPhpMN0NoDYKGulG/GT
fBrQDnuLf8qVWw6VKG57NSYCNncoHBU2KKzRdUe42nrY2omw4hbnbN/gf6Cwdd1g
KvTYrVVAyT8nTiibiurW2TVNfYdPDterk1SwMyBMnEnS0bfllsp0Gq4ys1B471Pk
30P6tXf6L1ioiKcbcN7OZyxeN6d3k83IkydvyUHxahBPZL/Yc6di7Zo398+HFlEh
MrvNnG8X5DT6ay43EGA9PpWyIzPUgr1IipcGrqJmsg3+dEYGr5E65Kx2R2Y+Nn93
O+7Q1kkh+NSCWHkGyxjWWHFNlGm/sykAnrpWK9Gku9L+gN5EexkVhOy8bh9xJ95A
xNR50AkD+Y/dysnPX2W9g7IuMiFBR9EMdWje8bnNewMsg8IMQV7skPkn+hw4Iyny
+QHtcnKuyS+yRA77fNkUH2T9zz0pDkRPKeSGzcMWEytnOGRaI95caWY6j8uD/vxW
QjuCFKu28e16JjSdKQbSgcmC/04RM9iP+Pw7prtCC/if8At0JfqE3ZkuZmdXvZO5
j/3AluU7ZejKadtV0iEUDLtd+t2mlzcbanvLcHULzRN/PmvJbI9sh+Bdx79BCkt0
Mof4ywN0vQgGfJm4v+QZIpGxn3cyr3OmRAun+0KKmMVi2P89n/dDyRa7L5DB90cy
KEoIQ2G7zQ1UgYi1cwGQXJXv1RrTGFTJ1TZL5ANLSX2EeSm4YmWtZ0UIygGE3pr/
fLbsh3OcZsnOXZrcgVEnsGMgfP/S2qK2AjLxTMzkzAOylIZ8OR5MK2BUWBx9Eg/4
TfeWNLmriZSLQZHhgGa4lp2hQohWkK59hbA0dK5Ptwa/Zi8Lo0Np0nX39ycDZ15y
1etDzJBRDgq60fkfna39+9UneJNNLRmNQrheYvB/ZaI5TXyDm6AMtvf2qBUlUxeg
fKvCRXqzk8MDZU3Qz3wkUer9DwgjDfwiIF3Wb1hsES5D8r2uynZdXG335/dJc18e
STO1EhGExpPkxtZER6dbB1sg9FXZ3rAH04wxA3OJ8ifuUYO6DAidQW5Gw2oH88s2
ZRmtlQjVGXbij9aBdwneNjd7bkG5cRqwfTNC4NsyhwFzUidgLcz982vXPH8pbeKA
s9AnWHY8AfZLi2uBn0/6j6pyf+dFNheInLCqyqVPeiPHI29pg9DNiNSt6Nzia2sL
ZggffOckNNvcYakoSlrgSTbXwwMogdix7mcpI4r2BwOrO70ws8QMZr7xDR7zHo6Q
XS0jKB0X4l3LlCmEApdbr4lCGHoAe7qU3JVJsTF0w7xZ8NnV8xhWE1aVGU/tt8Qm
jdGC3jAwGR7ZExf97rfyKOVjsj5uKxcVhAj2OffJ41ZAdg+A8FqJXFcGkXVFXvPx
`protect END_PROTECTED
