`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7x07QLZvzPiFlCnoRfExOTmsETSsdmvpzkukHclEBLKJVYZGPfJbJF6l1OSpi7LN
Jz2UxyIWGri8u3lU6QAZpgEhOOg2C92CUuNT0b4EETHssSCzjHbqrBir6q3FYnGJ
gy2m2lkuQIVp/4UR5HDY3Uw9pH82+HaV6aSFdIT72f0ZjqUHVXr4qeHox1OJiLGH
fqafkP/LZUzjnhlzhZxcknr9imM9ugbvbiBQAqfoNP8C2BCE3jj17wePXs1dCANp
his+yH8sD3PGHadkU2mszk7FYalGygUveKY/nkWBNhFIpEXpza8+VH8cdGUwbSd2
7u5qDelmgo/eUArQjIPH8uFZzXXfoTHp1lA94uU4ADpzrZMoT+ImABlXscu7UJ+6
dp1EzOziLIg6zyDWTXs5HS0an/htEd7T/yeM+UMFefMQCFxAT8c11+n6VuguOefu
1XynK/R83Zg3vHJQ5lAI4jf1tdelBP3aan+VuMppz+5SgLRiBNQhCtQNQmbkhtOO
nSE1Bc0cSaphOLpKq90QrqM22eBoobN/lpaD09NJkJXop4VK7DtcISJmFi4yhSl9
g42OzXeMsxHdTg+gsPznwQmEMVcDjO6kOfmIvuiOy/qh6JoZxB3g3jShMAbDJY1y
dbqvZ0/ApItdINQnuuW3K1K7Pt30DFFR4lctn86ybXCzQNrjxFt5IkaZMvqFPew8
lYVxrWSeZJmiUKyAz/lFK8J+qwdagdolAdaZt+XzAuXX6ViPmfwbMqQMU5MXWnQp
K2c+9xKWfsxoNlmNbOv6n2E1IpLXbTbLAtNzPXQ6+xBNo2rFh0IarNOq3TNt5YUR
EiZdM0O8ONSV99ECm5wEz9ZQJ8usU7bXkkODigYjpdNSyxXTouoOb05cluHpq174
prutxJpsQqai/V440khsMWiGoCkNNSHiqauf+M2l4mvohsI0gfou6pSA6/Y65BM2
TUtifUUeEuMmvPWfHNkhoiKRbyucOPTGk38T+H0uvTBUFSqNJ/eYagXV04rCgB5b
ERaya4AuRhSy+ktFLzOYYml0EPygD/qPMwVPH69l8PDJtbHdt3FZUI9ibSSp3wkV
IbjD0k0UCqVSdxPh6UfMKkvwW6jb1UH5xI3kBxtBfTEoqfxeuxui7zHJ2I6d8WXj
e9Lf0571EIotlNv3J9lqHi3pvDJA6qx3Xn4MDVmd376YsQNOTtri3VT/NWITX1aB
Q2I023iSzb11vLN3rDfzO8V2ZUAbNYS+iKEDT/xBQPn0EMt2dW0ClPJ9nYFP5l5w
1Gf/WbL99M6dLgKyL0mf5z7S0YmigQCxiwep5AA3/DWtm9H+p9Fhsj3KtVfZUIUK
ROcmTJLGER3GzDB/77pelA9UAUKGrPdKyvmuL6O2MvlG/aiEUIoTa2lXJo4sFs4h
HZwhDjNA0vPl7CaI4WkvwiGdl8pthqjYU71WC/m4JXu2ilVEUeeWOyalXqpXs9/X
hJTHHg7m2gltG2Jd9yVBf/PVkeyEcaHyXOqH9nIsoFStHBBUHIqPk08vOEBoH5Im
qTFA6YdzX6LEWLUPVZQH8xJ+gc3vzHYOd8+rH42M9ADTuEY7rYJ9G6WtSUD95n1m
Wls7tjiiMOYNhn4w9yfbA8z6PoiPz8PhjqAD/vg7mgTRkEs7zDAQ0xCwOkmRU62B
d7NqOXMH1oQgvFVPI+LH+MFEuEL8JwSgoICyfmBgPdsZpbKYut1nkE2LdLFWmQlk
jydWkUalYiGIaeHMp9c3zj0hWNXn3BBo2cGxOBQwA4zK+IzYcvAEvIZj9uaGzj5q
hvNUdwrs6205i4ceCNLvGLTbqTIoMnAIKeubaYzLcfaDkEszveLmeYx8evi418gp
Fesk9wNZRt+vhqEEuNcNl5tpg+WDAL8cxV+tandauyMFcLrgYvPlO64tNc549MUb
InaANXEePXuMH7ACic/AR5JeH8U73uU7+ufIaiLlQk+MkzGvoIqnOunv5xUYpaKo
8pV/tlj4IniUPC+pzrz2bqqpmyJLjBpVccvx9DA0YqzrpW0kMTj63RtC9wcoLBfx
CHdtB/FlI2/1QUeNIjP0TeJpmyaQxdMGqgyotd69qZXERcH8mMQaaLI2EkAyNPJt
MeqevQ2DijRK1RHo3NxSyiUPZhXhxTqWmbHVJ0Ta1Zsjb05ULx+eQM/p5GFTCgwT
8M/FUHR3JkIEsKv0x+zvHMFDbxB+94gS/b11+CS4X6J/Y+oNUzDYSMV+hPDFMt9G
g6jnxn7fJOsPmsLQ0hDXHw==
`protect END_PROTECTED
