`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EnyGYCcHHSkSDA7n/7vlgFcaZGH/D3s8cmL8zDm/0eDmmPhgTAUzRlc38Ag5fu9u
8+CMG9gSgFUzhVroBCKT8sFZdaHOZ6pN1UwinBEAmb8hFMyujODPmTUZTC3OQNGy
NQzjG5lEirwN6muFBZLm35lw/YqmZe8VnmJVx93/fBKHpUiQvq0XAcohCXjGORbh
W5PYhENYU968DB4gvGqWUz9CL4+9wUvOPh1O+gLZ8+O+gOacCaPgOzsIy9yaQoYi
xp34awCdWEP249qE5uyqpE5LnC0Xdj/mRnkIzW/yK2sHSpTOPS4+CRVoA2wno2Md
7EB1RLkTzcGgEEUL5taO0vSi1l1mdjgImvNBO7D5kfoOuVA6pb9HVCuSlxfNLZIH
GHcWUJmA/tqC730KTL6rNeN1B+3OPmlL1yCUzS9geT7BzO9Dx4MbxGjtYcRExFc4
OIn1P/dA0eahEpnHHot4ieFJ1ZphhKOmx+5qVEXI+XYBdc4LNzhQVOfYbMUiHuX4
1NM1wl+tQIBsoZrsdVS2/n813Owgtzg9hDkzWMjGBVnwDSFV17UbkPrB94NDs09H
zwYrYNjn2hmco7YtBkqhySYHx/9O70XhUGntkn2d6oxTLYRvHS9JpmIPO+21pTVH
oxAMZrUHud1B6BPM8Zeegw0IagSKe0MgQbMTCvIv0WuisZSjDr+ZRkQhvhepkHMC
7sZIOAXfXspACN7XmRUU40mUJ57h/38np3TzD39MNCZA3fWd0s5uuUrWJhC6hDz1
nh8OSmFw7O9Z4DWx8VO7Q50yExNGKoy+7/GCp9fgEPsXjNGZqWUHO6El3XC1tFUS
Nd1wUQicEMXjCHptyyt0lb94SV4gWoSRch4m3palepLUDWzHERbhraYaYNLGnKHt
plkYWA2iKxzBmT2YIwS3YzXpdV179qy6sm/FwXF5BIb4XLdDI34QaUFYIOmaatcb
LvoCdNQBrJceSoPmAmwqLClUEAtbPbKZGLSt6tze6Z1nNMYtZKBVLk8Y71Zq/PbE
F3kQd1Wtt+gR/xhTMRmQUvXBw4Y3QAQ5KSlRnCtjpZkaAWbhpaHkd1VLL9galOCz
R1s0GMRaToDkenaKSO8KIf//f8yXcIdpHRxIWhuBca88TrET2fcvVlEdzkzPZRUi
idJ2PemFlvFXYIiIIjozjJdL9RrSa6sarQRs4d5iciFBzD9RW0lLqKHvFSGESWBd
LiwxiBtw+d32TLA2/8T/DNZh+LIJgiF62+OJ4OUht+8I9CHYMunbsTD1fWMDd+21
mFk3inpbTx30/rNVHdnUVC5IItlwrenco6rFq2ZX9dr3v6tYatX+gf50C8sdKGkw
J6xOqBZM5taCDR5/fMuhRU2sOCgIhqN2sIlMHU729W5MKsdUs+dgimIhjFKI+Xzp
4Uw4Cx7IVLr+PYvMzx83vWouQoFIc8xhi9/UoxVKnaJXHb9DQigBRhoKnwQ3JBUw
7cOxgqZBQNn2QXJ71BkIMUGQKrDK4EcEkWzxTzh0Z68ar7qarJUYWPTGQDw5yqJX
YswapaegovTnanPcMa59ii5YOXeCJSx2kVbpWTI0oVT8IvZ4GqHXeQXAU+s0R1K6
UnA0XQY2BFpxhgLuDkfHnTZkyoEZPGO61738g441Ye5QceC72LwlYnw4/wR1YMfo
OZR6L8N66Sge/sTeipS9MdlxkZ/fACIx7Cn4MqWKVzU/I/2vzy/+d+3yOMrMZHki
BH3ie0/rCDOUbdh8k20TjE8x6z4P7MmKZR0pV0QDADBdllVYtcnxFQZPrCZggWDx
dLlGm1rxVfb/+gkV1Cx/9dxfJ2LLYf1ZhUsSG7BlB0fRXSW5MqhqBoy0rk1Y0Jsp
dZcUcucyQMDsDLZ7xiKYPEzhMNv4Vs8TBvm6G86IGvjXdr0An+wdWPK0GGVqJpau
MWLpzg43Pw8Q3SrV28YzCaDPKVug5Zvso/g0fvNETYnCpEBR0cs2n/KXRvoYCxdW
N/FpLv4Vd+/bH07YZSnYueom7ACnZUx2aZ83YAv1QD/iSfkaOTC0l00mrq4uRcgJ
FBtqA75VoXO+WSxuwN+v34Ysd4Q5HrjcT/6AL9JO1LGB9CJ/5Gio8iDevDVAJmFV
opL4ohl9naAQsJ8aub2fAPFm6ZVSSs29+9hjKCUuOt2Xqd0mdX9btx56n7WAsZ9c
c7qWbtST2dI2OiEUBf+I5WoEQLdV7Kh4KKCvwjGu/nr9xsgK2e45hEO4rtr1lZ0L
hnL8a6U54m+Qc74doNU3Hy0ecVe0cuhblJIxCnYJuJbngtTPV2SDeGah4cSo7bbQ
jnjkYuXdojNzeUoTcFtzZQTLfKUBYb+4MbkSOazr9TWuGa0wE3HUoyz+OmbGGBEN
b9fpJEjlauwZAq/URCfdkNix9dtv720PO3dNAsJD5TL/PsKE+OEBbU6ojWeQHZHH
dABVlHR+rmnyMKsCY2+attRKBlgTVCFjWEUj8IO0DjAiyMvpX2aKEN8Bqc/ahTAG
7yz8n5h/melMwuzOnXfD/abTxx8Jj01lS51kmQuCHzYe7ZgJpsc4fHQ4mY3NENPq
MUdXNT7Qi87+6E108Yfp9fvAD9tk93t/MlNa+X6eAx01AQ+qVy8j8//nN/iLRt1z
JL+v8+lvsoS1RS/FlFZUyWnH0/H9SNl0D0tZx7maq3bHO9zXT1VW+vMoHumYSNdL
UK7dkGQEhB50hrARDm9Cty7ov3PUHNRgROjKVwC0XePS7RvhQ1lI/ioHEuDc3Ci8
kNAVYMBoNatGpQBraa3oKobfA/t1oC3813ORgE5fTVQuA6u5/SPM+3V6t86MnORv
Rqha5ix5A0m8NoJKgsMPGzdS2nK2gHdYvmko3C3RcZxplY8zRMdYFa/PxnNESysT
Hmh4SmVfHd74iB/uoBfWz5CbmC+IGnpTuW4SXfnf7WUhfTXthaMFRe7T4L8/6/GQ
zesAsgZ4DBaFel2y3V6Q3QMPbPA4Oh+eBV17IlalLrqpIdk899nLHvp/VQ8RAyDM
ijwcAr5Po/xMVDtUD1hYxeGSBCDOB1iiDmTijMFSKdcuXZjHtErb+vLyFEtZ10tt
yzPeGyFp/Sw0Jaa6+0+OMHM3qBG8r1rIwtnuT1Q57gDokG7J4dMnNphvGTh2/RGc
NpToUQ4i1F0p+RQ7N1bMB75C4IdwAKkcLUVRuaDkBlhpZKkmO/4OatiFFg90VCct
cItVOwGizC+a0WLq2M7HuEfV4S5v0hUin5/HIf0unw96pnorK6uFJ6+Mhx4piiHs
jdUiFhvJl1fPYVYKDCYLfye3OLLJyIOYwMxd3o+5s0Omh8C/+sOtQcvPYTOdyOZ6
+JlbTlljcwb2fqZX2b4Uv3AkZeiNbOdNLByKdcrCQHcfb7V1P1hz+21eW3cU1juW
cvoGZgwMrQwPoPBXf8/8JLitV/E76LNYdGMMvBV3kjmfYuFEqDzrJkrrUwlooRcG
d3Tjlc4CfF6PSMhLUVcHmBJAUNDkhtQnHFVZCNWmslUrne4bnNlMpKuzfwlAFdC/
WVS0I1uDuVj5pJDBsZ7qYyKp58ICADrk2ESZguzQB1MoZMsPhwVnDdO5zXbF/MxK
xYbWtV2+fx5LNoj7MLQwUtV7lqj248jlIUFxWMjH8/gq+uA65DBJNCsiiCodT5X5
+fdsngxnRgY9hcPGf3UEwH2O6sOs2mlrVNzknc6HNkvxneCqi2iDH8XX2aoWvUR8
Dka1pU+Ie9tbrCfVnjpl5GxC0OZ4V6n23ZRTO0uK4F/+q7c+Y3kT6M5blpWZnPFS
BURgnOL0sDhXdW5gaUALb/Z9pamoUq9Wn1bUIUTKaz4CXXoeCkWcVCuQUySsFfbX
aTkj2QyljIfWEHN5ckD3sFZd5jhZrgLUrJPWub8uAhs/2WGwEiQsou+OTj7XI1Hw
1RsO5ZTZ2IFMllNWSswCP7eRcSLDs7g45rRYz5l5li8A4T0UDGtBbHbMuBkkYZhM
/Ddy1KBED4jl8K7Wmy/B7/uhkGGuwOEeob7IzSM560yaHHbPfSfwSFsGbHYZrHIr
gSrUZHsi/olP0RVHFtaLDlgjdn5W6SZGu8YfFy5lcz08ARoe0gATjvP5QPUO4J6m
vaF7RddchQKXR668SNiniGPKL2GANcdZjP1NuGL/E26mvMWa13EbrveDcfD8myFK
HqdM/+OIJfHCnKhhrhnsy/6KPQZOyx0lIbo/NXyz1r9CKPW6fwohps+4duEh5tG4
xO0/WF1Xr81Gzo90fjPJC43ABKVtkfG/t2R2guN70xgfTbJv2Qym0PfQJLwYPu8g
LYt01+SasDG0SLrA+/qBc3JvvVK1IKgR3M5adsFHvmef9fYbm87vGvts5zW3LVvD
7z4R5FQBSzQFmyV4819Jdkl1+ks6tF24TTwiFO2t7hL9UiGXP+c10FjVPUB2QyDk
XNOyLpJBTu/0NR4GUsasSF0VlmwCPAVJOTegEXcuRJYruYCnF5KcGyUuvVkTgtrU
0a3JMRmwuBcb8HlCOyHMR5b26nFNHp2jgjJBUyp9oogl5DD5hiUarc0Tvuy0g5F0
OpSPczmRs2GZyHlhuOlp3TxbQciXuMGH5c9nb5+URmmpS6iqERtK3CTXXvpZCBm7
lucQEyyxrM3psWOn9giKEvZo7KnTvpFMcakDHtVnn99Ekc2czpGsR2Fl0+I7NBk/
5ND/Xuje+nVAF913dDV2hcnPzS6rMqE6kDw4rBvxOatX5AalbOO63WxqLqTeu4QJ
dJRfpKIvODF5Kw0wxBlEeFdm25KTbA40LQ/X3dsMLE6NWxjHhFTs9MRdV3Nu2lLZ
IYnEcAbcZG+Rd4ruco5w7jP5x2EU24+V3aklEbKftBTcdocopN7yYl0hKqYZAXL2
Q/CPUvPhasliFuy8dL7NmEAUvVUHxY2McZRaGbqllS8kqnRq2yimLZwUOmdYV4K4
BIpktzF38/2bUri+iF0HRhWmm7XDV7UgykE7RLmWjrPjNgwSDjHi0i17IxkNZS5y
a2bnWpQSM4gYIFew1UwjQcSwlv70rR0R18uQicKGlcwrCBahHpN1d/ffMqILz3AL
6vuU4L0vYoIvko0UZujMFciPup7XtnOXFoP2s3Z63w7jK7eEjGTslPrW2zJur1AR
n1jx4bNJ5tTeObQJ0578oQr8oEC/QP1CLUVaS2zVzLnlgLqZolYDBMun8FTDRdER
/JoTe/chaeXbdO724njsH03pRLnSMAAWhtrz35JZbmrBJW8Zqn69WdHYC4eawZxs
P7SCcP/HC0M+HLlHRX4fsVimu9vyIGcaPNLmILoPsI0ZauEwbQftXYzmeYPH/Ps3
eI+ZBnKuBHJbeg0rQWlH8FUXIQg7CX8njeZfcRa49ImhPhVacWJPYvWd9XEllmN5
pW9/XFoXyNwzlvmrxo3CMtLT5YJRDwx7vQcRXbScyT/9NPHzpIW2wT34I0pnt06V
HyLEx60bzSje6Ifr8oA6kEeyf6MFB6AtvyJKLtvvW7zmAL+5dFaNNUcfaVdgnzN+
CbQYk3InY2AeR9jyNPxA1x5de3pqArQaVmHuUnUdeYvSIxe/LYR+En0lVcX7bEI6
DBgShvaSJ0mJeGJniNKqamBe6cFb5pRS6zGLXGbz0Iwk6VO3AueBiIwWgN1OCnsg
6+20b+L7QjXn+n619LUVW/WHoSjcnchx5iwt//s4bqlxI0GUppNkNUtcW4LT6vVK
iv3Uf2izcosf52XSsZyeZOtjGQ86iL9ZSpv9Qt65wyUrUaQhgKedXpfScyNpZ2fJ
cnKrZLhS+TjgcjbWmy2iybhx9R7SzKKCTZWc5ePHvRihy09PV/H+wF+GSmnK5oYR
ndj2KHHpUpOhkrXOip2qjGFtvKdoZ3EVpP31xJuFCV9qVc7r0pdqE4oHk6AIXrmX
EKPy+h2QLIEVluzyz5TNSPtAue4J103naJ08mumyS5EwJrCswwxSg+QeJ+UzxkuK
gC4Rnhyl1cX6TGrChIzu0vhdVjr1JeWx7VrYv35+lDz51GPW2BfxH1hqPHNYlBXE
BauHLIn6yWdmYJZyC77lMIvoO4hZRNgCS171QH5mvM/Co74dnWKk1PY2dZ3/YUkM
z1ovOCFHDH28Mnufcx8yUt7I32R6PUTr0qx03w7GOL8hWRMXrQDIPWNkGFbpIjnK
xfNjs0hqOYlVqA2CQQdwAVNVhf9U9eosl7zFL8G6we08ZuR1FM3rA5UsuMykQCxz
WR0ngW9Z9PDUYBChWIkA5QRECcko8FWaHGUb3w0gzKWZBD8e/6IzfyaUY3fhPo0l
fHao7gvRjfn9xJU7gbtl8ew1kgJ5fJ0yMWCxSSlAfHKbu3+UrZnykAUZrQH1bkhp
zdeqSCUZC2ag7dT0nvofVpyJDW9mTq92CKGkQ3f0hqY03z41dAYfDTrVgyhalhwm
K7U905kgfT1m2Oh/iLSCpz1EAHqc7rqZxJRdRzAnWn+AIPFvPGQ6MFIAmBUX45BS
dhsldeBOXN5L5u9q3tFFvrR+1uetVyPxInynYzyjl6I1cQUqQKg9vDJ/e8v2Ubxz
s8s5cbFYmShMCj0HEmND94uPOZd3NEV3R+mb+qWue18nrObFsxzY3hCa6guPtgcL
xYHwbqIrpNn6aTUhlU12XAdRQ9vhAH6MgCUQC4B3x/dPVfVhBSCagdzIZsNEWdQP
hK23CEEgY+zDzqMfIceWG3IuVkv23n5QXtph4tjK2hM=
`protect END_PROTECTED
