`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JF6hLGIjfO14+iQLgvVhE02J5VA3uqqOh/HHowtasZs47Dekt9NHnqxhMXy2p9ww
Gegh/dDiJnI6pOvi9DZDMBEoz8AFn69LcN0ww8gD9MA7g/pMUEkf/nNYPXpZPmTW
WxBP1Qm0rDF6QAlbonMSWZ4K9TtiZrXCSTR8COsxOcSnyxzlviyWIIE401Uxn85s
AvZpYLTy1Us8/fwqNq/buvmPnjIHmNzsUPXa8Uc3PUFiOxq0geypTk0P+lzoVZ/1
3/WaSRWB9TBItXYRQ8+0U87yrve6uULEs/APuqrTwk5uaqqA3IeanhzwR+RAW1ww
dtjpH2skNflJGVmEOM/ljYtSxh0KeYmb7QaeF5UmXmwxxXd3srIgTPZ+NT7eroaP
mQSSxSUcNGvlt4tfF6iCini6RKWdRzMWajvv9rjBMCBeDcPwaExBWJs4Gv9R3z2c
LZNsiNMCFOhyPaRFsN8EHM/cUtYCMeKsr4OC4Y3AWwCRpTkXtPa2igoXz9l6q572
KPK8t5NnusAaWHr2ddbHGL0MYg0vJOixalnwUxUg6lU764G82paIcpTqG+uxnOIT
g5nBKtrCQ7l8NSzFioV7ePfw2d7Z52tESIDj0IszBaHjT34Dz9Nu5V/E1eJLydA/
tb44AYa212xH4lfAgM12PV1Mr4royj5sEm3A0aQd2jmdHa2fJHhvzDcULwb+5u9D
YLVzNWcjnz6MzIp/+xnWPmvxo/n57cFKJLo7QWkYAvmzDI2Pof9j+cJwa0ClXbrO
nLy+/3KrPQGvE4Bx49s+2G3vpYY8cr+Xif0ip/SrFBq8hpDPrTjDmLr22W6t7abE
W6vDg3ujReGUyKbjKu+rSXS/7s+XTpjfhEKbkDEhJp2/oOPNlS6wueMrtNHwzmAS
mM52iLExOW5DPqj2IFw7ZjcB7UXWIyPXQxsa4KcMNdgF9ja9IUGW2Ns70lmaZ9Ko
nqmNuSQmQoMjhp+AtUSlgxkD5CkSHh5lyLH/jcyYhx9VriIS3grpcduG89srHo5L
hIHA9Or1ZsR8ive4tTW8sRZLw5xAC738bA8RIWvgV7hY3C9Fpe9AsruN/GdVcI4P
SPlkxSTUjxWoFAqtUls7Ijg3uQYtnB/vB6nHDapZo/9nq0GQ5P2N7Y2QWHnFC4VJ
+UYpRCQhSystAFcr6srieEEAYJcjaIO8L6Xu04tGzpDloztFK8BBcxtTURLMG1dj
vUk3Whas4OSeoALq4ffK9buWrrnG1s4pAL55c4Qnhzbwlmct/MC6fgXxGk0QeLij
UXsiT83tjDBhl2fV3b/dNJ3MvKMSn/QkWUlHqHQ0GpATysbOtyVFeTuzOs0qtT3G
F7AOYrMochhXnqcQqFNYruu0dnSoNYYRArcml8mtok3gJJXS1YE6+u53/2kKAFv0
jLmE3hM9Q8CFJAmmaKF52O10Yg1LRYyZqUWpm3+UO77w6OdPeC8NON1Se4opppz8
y8q7wuzKSOWXhAEJmdS+oJJ3J5rP5pxfBaWsG39wQ/NwEH1v9d8LMF4FViigw60j
a0u7YkPun0g5e9DZCFW114srOGGwF0CEMIhNKAWRTfwDK2piuX6aVC22RVnASwwj
QpZlMRyGvWpJw+FkxFk9zZnKb7LQzbtLzrkUiEseXjrd7T8Pho3fpFZCH7zaF9rx
hPF5WZ+jmZxdvr9kqsy6ob1sE6o2Q4bF+db7K6jmYGLU2Ae7Bj69AnbqgNX5dHpn
kw2iwCPh2HHX8hwkbMI4z7jICD+q27+cVqxBq1IU8my0y3w/BUg5fUgYqMZj0RMJ
H97GR9BGpOZwIDfuOy2/n1i667HpEuJH2KLZCCUBI8/4kwHM7lV2aCiSrLwtbWv5
IYQF6YliXAeIhpxdAYwZyZ2SK5lDvkz+2UjGVZP0VLYhZgmnESvxkbU5BPxT41eC
TGuMgE79tY1lNseJBMV3JVFF7JLSBxX1Y5DdmpNyU+h1bGGrdPg6P/ZSGc0al47f
/MnvT8BuJOSPQBy4At1HjkCfGNZc2zSZTuwq4aFn5giK0gznow1iUBn+d87LsXcH
`protect END_PROTECTED
