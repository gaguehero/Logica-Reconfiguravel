`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dTdIuTlDMG0/wrQ7yjEKOlSYzhDGbfjmP7L74aCpAVYGJNsx/hlaYetQUC7P7oZf
A3mBm2BK2wbduxEy54O85TU31f4pPCMEO+gQO3yvafMT1U3o9XhL44q9pkChCuEf
3ucW/P241YtN03Wj6GO5HGdtA/dsFcmMroiE0nVl+r3V8degn+MXY5OA89vWpMrs
C/xK4HA5IPzHlfVecPNuBl+ezV+StDq1iq77IfVzoalRCdk12/5aG8LQpXZ9O7z/
zprNu4BoFqH47hJSJuILKvN1WrfFoJMjVVN/OzgUYiyis76VWb3kVEhzpRDO8cAl
UtDh9NL9PL+RhhaKaL8cI6IFOCeKOVSFU2q+vD33POmWzBCdir4UaQBjkP13bzNJ
qxm2eQu/LtzhUnpxKWYRXeKLMDrcJ1PVunrXyOH4Dh3PQiew+6STST0yNuOge1LL
8dW7HFe8lR+kjOxI46yAQXC/902I+ermQgCDyz5b8XzTvb7/dQE3UgQX8MbST/Jw
WouUDl9Q6/P3AsUMFqxfpdb20pD4c6CoeZsdny5a8UYyXRd383T3Y/rewicnJDx1
sufHM5iZfZwfu7IH+F5ZNlqCp7aEd9vRtqUFG4ollxYCZcnu06UEpi76xsLhrFnV
vfQo/QGNbz5NR2xYYDvzrtZ+jCzigZYS9ku99JFlV5rOBuMCp4XGlbUJpCcXcNNh
XypolZAK/VY8nb08jtPJDwHwEgjJJVEcmkbn796b77rSnlJH6wP3UFkwIo/zC1W9
5V2oB3x1pUaglffXurQIKzl5IyOihBX29uNWVtgGgXRQH+jv4JcvdrLxj3kny2mM
jMoNYZIyYuokmxIbtLhG28GIjKNElutEWO0tgTcCMWDBYpNggZ3lgLRPpVK21mnO
y7vQhkvHUErOI/LIVxkgQ7XZfF5acL3nPqA0lzE9GJFZgWGsaGADzLGinXfw8qL3
7nx6Efwh20Syg3naY/5BY0ETzRa5QqyKoZ28T8I7wZUdsvMxLjHLuIgRxvMVX8QV
MQPCGQaWPxLe2kgE25+T9KXokiPow3RDgoolYPRwQd1CvzFIVZyxGHToIuBKI2A/
0QJwEnD7npmCD1zI3Xx+iiJvPmusSP1gtCHO5Wryz44MN5yezEnha8gcQ1/dZdvh
IWAvgEh4D071r7cdjK5SPdS4uI4qGRMRfxIcQX5Q16aQ6/AUr/22WtUHXeGr82Le
9wo1KnsS1Hg+LLNInPi+qfxumxLNkPpFkLqbYqEaPjRpiOifVM66Z6xQL2WBJ2Ji
BUd/mTrzgBalgxSimzw79YlF7ndjnlLkqQua3HiNHf4QjtJeDAevFeQBXcoMV7uk
Odt4YSWWXyyi7Wxio4h497eHOgODLh2Y5Y0GcAwT6QWeGfwn5VQh2O9jgp1mdV86
yvSWNDHySKMr85gy1NsDWzcKFOrVkdVXS3PEMJ396fdi2BLbW1ULyEbM1RHaHqyN
MuO2tNKF2PXrgru6CdWxmYZpBDcRq8c6yd24jIGoziPxGcD6AWxwblCBq7sNt0Vo
Ad4ctffbok+LafWiO+iuv1NbzntF/CD+CUUFIqv+sTvQ9i8fFSh9VudSUSZxcG5p
pPznOmDI3qJxgrQGvuSDmH7rdKjzIcm0qM0qbfhHjEIMi0TCYr2v6wpoV3KUTOxV
SLbEkgnBKou1sSp8sVJ3PkPaDkafc+l2tJZpaw8spnx8DpovCtSpKbH6rSv1REuA
WFHIVj48OLTPQJ8GY2PaZXvQ4VzaGzq+mu88kmpj3YJ+8NrdATXlUhGYE0Do1kU1
guNC52Q0uPLn/9vQNhpAaF8ACm8MFz6RiLjK0O7SsCtVG/9Y8telKDlAoGh66yah
HWB2y9jTSeHOb0S5WIzsq7sYWZYnwZo65Jyh46Eae/SY7C9Q/6MCgT+CMYk7nnKp
cyTaiZiNaEFhAteD7ODRuwkAVxGNGmuJnJaeegKZv7Q1rJilvo1FjDYVXWzQ/Zpb
FHPxgM4s3xvPmTQsR5ziU9Hhwws5Oe7H+wuftOYFUkgJtuetZStj2eTL4jubeB5e
UuuzlK+EGjASeWg1WuUkf8FMLEmwlZDPMTLh+sk4cjNO4F5Eon+DztbRKNPwSu3L
XKOHjS3+gaxCoP2+4p9bdfFtinXgpkVUw22xlDKY54kzsE/2EZla7mkR4MhwMU+Z
q7kWPu42nEB8zKZHAiUM34b/YIN5gz+cP+4qmS2qDi2JordVorYudfMp6j0OFnoY
wgI18eV/KCR8pOWBqCLy5rc+wSFhEAa2Zbg1WJ5zB9zX9l884pgxACKRGMrIw1IQ
VfE0RkEqH22aZRcCUXdBQC5KPwpHEq2rFLt4hamxbGsIQ1tQLBb18/lA5aCOiNvQ
xkuAotYwddaRmplqALHEyYequjUL+kaZmb++LgvkYJzsktcJLgE32WZHvfY7bAT0
axrGbvdzGMRU/v64GP9F+J5u/6W+nt1x4HWfbCSetfawYRPjqsxGzPcBaBtgOe6m
F9jPGb6Mwbt37Rgxe1JZVceHEijD3X4WcNpR9YkqR4fs9DBx34KYIHy+BHq7Fs+p
3sPWfkIcMhFWIyvJADu/swOv61ex5Jas5sZ21LJEsn2wF/sLjFd3ba8DySp7RBuB
T/Bk8ZXBCSxm6mzYjVACQH1vbqnYu/WuVsLV09TLTQmESjHwEsQ+mudFpd34W1N+
zSop0iJi5omAg1TKBLGMNlWwL8/paMcgo6XciDyokhRU1jILebhNujRs7U2hSEKN
f7jArESb2urpBP6JbQ2QNy3Qp0zZ5hYtN5cq6+BWSdcvizm88El/QlMGNJcjhmmF
xrHo9n1CSPA+rUtNf4svtuSQtT+LDcazJwtSF4dnhldtHBYc981SbdnLYsEUurJy
fCLALNC3m8mOxVS2LC8YdMcKoqCovXTC90lRbtS1WkrDcotSp28mOHOgME5XRNXC
aciyfA6l1tfnDUChj9XpnB2HyjEONiwcYa48VZJJQB+RuDJSFcwMIPGjYnXqBmz8
neWWvPUogBfwXP+0pICJNgZx366as9AP30d2/tlUuUcyNqP8UY2dAYQXO8lKqSMi
8kFiO+MhkkiedZBywwfjm1r959Qf1P3lA0bv8otb9mCVfIHcWkJLTYqXRLbKHvEC
/Ebir6tQQyPn//VPHRHKN2eoaOABj2gPyLOaqwZSxw6CZ+AmphgcQaVYl/9dx0ZM
P/QKwoU0ol6XVAkJpOkpqUFvWJ+CBmRpHCRrY3VkgoVnt9hIrItaHTTtEtNltVom
6aweQUtta5LawTyMEq5dl0C7/ByBJAXO9oeX37FRFwEe0/+3PS1OBJr9q6gSe9iC
0wVNEMyhp5TZLvJbXfIeWNPWHN/w4MnDybdRlTXIb6moan1r1SKnLV3dnP9oN3Wr
W9QnlLPe1SM/E5DCE52IpMMF4H18479S+kzLtQdj67gKDr+5KU0BsHo6QLcSEsTc
sapPGt1G5/LhI0LefpfwlrOLT4a2V92o8POM0LcFMfwLFvfNCrZfKiToR5FlDYvC
b6lBE6bx9WaG3Y5X2qxhEntZ57xB4HKuFAoWnILNEKaf0F0M6Ja/tRum6TyemFmS
2cxOygpHwpQ+Nnoxrq8RpYJ6RZA4oSsd8Isx6A9ZrVnZOxuscyf1VPi6jYlwvhPU
+gsdgnMuD8wPWxHzJmGfHsHxB1sOOyUaZSmLE9JFYRgqgYlUpvREJScLclGM8HvR
gtb6B55riIrOiFgiwjYwbCKdgRh98YGpje56+5/pw+aQubtFIWOjQLROPHlobWxl
u0ggOmCObZXeO00i3GukORl/p8yRpOdbYkg3FXJRzzaA+cShhFDR+VvRVmkKUvfk
vcNKYEHEn/u7NzW+GNlCkSr95wVlKr810UVQOtLLjgSBJdIdVG3MCxZEVla53y2V
mgzy+L37nER9dJnXsLHA1/HMBN9THionTHf6gFL32Q6yICvfHdTxtKaL3wcAfAhY
bd5A4vA0WRXZn7q5kB4WmJbEVZRycGuQua1k96pAFf9VpNu66j5V0/JWjgHL1d03
lKqI8KUzvXCYXoNeUt8BIzuMa3ZHu859o+0at35vsnEKUzMt+/0BR4U7h0p2Fz8l
be52ZIa5F/LKkuRq2F38LEjqB9EmfGyidUPQm4plsj+Eb6s8FkZKZ4RrAgBLu9A4
K0MKVSJaQIpd7htuOlcBsjUN75jkKRA32D3LI8DAfSTfC0Axj3JXw+tFu3U0mGQS
ZYjrGhvcpylFpLAl2Gt/odHqsfqZb4WXGShzet8SKcwYtikYxOJgXSvLhvcXakQZ
i2vke+X4NMtMKagwbstJsqm8mdIfw647pT5GELnh6tvPptAaD3gvzB2ycdbrcdL4
b+sg+CTv9yq6e1jYFlay5Xu7jT/zjqLf2qrCb2+NUp4DjhhEYGhe1k0JSe9TdohI
ZA/ympOKzxSD7/ChbvFwesVjvL29fQXfC+5fAEaUPXf4k4i+sqcWuiu7vMOZVjCw
NUOqAJq0PlIT1wt7875bq52ecDSKjwIvlkwqBObFPC17Re4mqvMbPP3t5869mR+m
XbXYMOb5LiQjy2PZ/GCGfzzvdcCwoLVtG+fRqzTtvJFwW9ew2nNDlwgHMRz1d4gB
H2D4HsuU9SIrb+niOLi6/FhHXc2xc1e2zMpLroijxSCDZIJfZzZkcHEQjwvxhxrZ
ViA/o2VjQvvDlGmvkda0FMmtmGT5lCfMV11Sg1axP2VTWwe1rpmdRSAnEd5YjGhj
Xkysxr0EN9zHVjbvMUKvGWUfBXc8o0Mn7rkJpFIXqrM4SrEe4z3nwE9uTDGAGamL
JHGkLHNh0v7O55FgllQUtSbQ6PShRhgX0gFI9NB0tq40MId+GPIBqc8Ebuy7L5KV
87fEKncsbR1qdGRSHS+Iv8A6tsQmMLrpMFM7O2MCNClJijz5qm2Nllf6PnBxVekR
/t4UyIQsxlcL7TQ5Gt2VaU0878zOkyVLR+kLOf2s1lCW+7epXwOoQsXqMc0gorq/
A5V7CLxWCYd8BIpUTToMqo58Lo/Lg0pEURxb5NURTQxNjw71pXvixznbrljAS8D1
1i/RlxnZP/jGgxC3ZFnv5KKr/GTWPoF4smzfG2Z5u6i8i9QxvuXHdy0WRf2/k++d
dzpr6tkRUgVXm22mlVoyZIw7toTYcSO6hcWllLlv4gMsJz4ds420E0A1/7Pm/YTN
znlAAq186wKhEvbz6dxp0rYtSqrJDTFqUEF+wCTnPGJ3uxNR+DO0aJufo9i1dBcl
5bl/E+DX1u+AquEn4ld+l8hkzLjDu9CWa4LE63DO9WSmL3xfuJVceA5jhGRSDyKI
LBKdw2sj6gv+lgtqJGLqYi+dKOnaPhS4lQw1b6cQgh9zeNII4plv+Ct+BHGlrZPx
FeLpGmKeTo0y3SMzr5uwsczEveieVm53eBoZZ73/B/Y+5MjqUgPC6p5IG+bQgSAM
U+pzcQ4pKty2HKvocTofz5Z6oknvo3vQ8eg9+nwJLbKly9hMYMXlF3RBsyNKbOSy
ZdR5xZm+fp8aqerCyObWp8FhZzaM62xTy9wY+DNYHHJtuKbQ+ytqyRDmc1WaG4ei
qDGZTRgptRC9d1sW+5eaKnhP88O2UupTd0Om/AaQI7YYGrJk275VZKS9W2oEhLAM
FZyP52N1G4oYSK1NG/FfkXeHxfLku4vEQhSnguXpSNPx0lmMq0stHA2cxtR2TQhV
`protect END_PROTECTED
