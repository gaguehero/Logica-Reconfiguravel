`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVXuuP58wEISlHUVnbhXHqZXPeqBXfBNtnw6vGdjECi8Jmh05nwns1F/VZHQXkp7
EUi702NMzRq96FPFn0hJ7KA0yyHsjf7zG+78Jobx9PuvB61g9xn+3KV1HPxZA9R+
rfjTHXhgRbW/KerYoxUhYh33e1qjdA+NOWFPkcgLSQSEwckkMqEun7tsgMIdWSik
l6fcy7P04sg2Oi0hcj7siMg4Ch43Rjfj4PKJos/ErmCmELZRFWKxYK59Tf2Nb1F1
Af+YrQ/f6vrkzUcAYhhzs1R4smJ85OoBVtwmzbTnWiWdm1pnJe4OwCGRyWLFYEkx
xQ+xmOpzL73i0ggHnrj1VlmZcVw+BT47bBDEXLQTohFjFj2UkAeFVtKZ0akcta95
orjv2KA1eSxZDlnfyytcNvc4haO/GzkXxfZyDoPKtAA4EoJlKmZBpaUGZfMmCap8
XhAgMPFBI+G1k+YTn5EhlTl2QpjSHCDcz+1P+Se+8fRHwDOiNaQnjby7Nfgs542F
ZaL7NlAzOLXOth5GcoEi9hWrzMpUWP3S4BCWpsaqjfNn0wlDc5cGA963Ipi3/gl8
Iwu6Mh20vJD7Uz/v8vM2TJ3/qjLHcksZUg5C7W0a1vISPGw2dDKs8KKWPnGW1QxI
3owc3YTsi6TlsqTEveznRF7u1+7M/OQfmSw3BXY4/jxd+vkek6PEAw/b9PX1D7iu
8dzUUDi04uBmYi/bvGz8mqAUglUYbKzC0/MVhQNGLglSB6iFxE/VK17YOPJqQfUG
mbuNwrmW5hVcWbZUkf/WBQlsFueWZEX4nsyaDi912m46fR2CEITpBwd5eOBxZwya
nMEL/v9M0OTTWSj+Amtq1eRS8lIqDdA+Wwz4ChfgogbanErNaN7SGoxzGWs1nd9A
bh4puQg1GcnRpN8gQ7hCcOrW+tPSHoUdD6XVoO9DXkI+pyeifV1alwBgqn/mYM9W
q8ldqHI+CX4ERwWw+ygR1RP6yHpucfuc+4NgfRgFjf/C94e9SL/d4UqLHDk3GBec
kSagi7hfe65CFWr70OMz+p/Nq66bdrSrhyT57p3NMCG7/IsTTFw5NGXjXnKKYvJd
plimWPiyBZ+1gHmXZQBzFHfou+FDgg+wiOzKcCbxgYAQn/GinNYUMKOG8j6e3u3P
98/ApebDV+Ns2hdsFIZecqiFkEG44eX1ttichEKaUcu6eWrVo2FKpFp0s/bnQPqL
KtZKMV7Ozp1Lzs505shHy/9+p8P3UizMeuekbwEWaaYgmiKBtOqD2725sqPSWMnw
ee8cPWvUOJpjOhbEMre4i9F1+cx0VIEhAYTBy1r3M4xjq5g++TCr95IbRwGC219T
LPc59ei3OkJW8aCCrkNv3Tx6Q2l9XVrHaYjVmFaieiVq430D5+ZSBpUJLduUC1Wm
TcI+gljZRx/c92H7oGZ+rtz7Sc+5zzgvWQk7xPp09/2NUt3nqedx1XoBU65rHOUO
4JdQixEoOhVqrand8QYKgOdAsPQA45G2JrFnoUpsc33jZ4BluC8DgQwAST9ZD8n6
sje8a0Rk8MmqncivKFt5gCJS4gJwo5vYv4D9LiD6Y6NZ9+EpS5ni7XJsXlwm5cEG
wWX01Kq99mtNOrCoGmOw0EScxapmPbLWj/yWj64oDJEOR6tFAMKSI1st2fUNUsaR
+X74K7j0aNPx+UtnfOzEn+3dqcUJKJM49MUBrTDwkKVHxrWtvrbMBFQsaKgYj8Zk
/R65DQaxElv74pPKB/uLyrNbQWgRnujaxMGkSmMMlHM9xVulc5hxwaTW7cvl+/d0
+VkXvu1J3rTODTV0tp6f3h6eIuUXS5soj5zuitVrKwjF9QNRW1gDUJEcTtxEg77F
zfdWAFWf60SQrbzns4D7XPClVxQeF0D/+biP0OwtPV2+1dzOp1iKoON6XQ52Onhf
+Nf61Ul6aQHC/L04gfxu1HuBz6fnr65ztcbOpyqbruVL4OP2OjgXGsMI9GiVXqwz
u0tsPhucDbEvBeMcW6TukXYiMZqIQbz7isiBMqEIPh3szvXlYWaaMLdWEsH9k684
19AJrOvdtnlySiK+V6LEqGdocHwm5yQ3i+1okeR/0tgT8phShk1AHDP/OjyfJO+P
KlCrUzrKYlGnH9gWlev5Qij0VDNZSxtzVLQUX7NF2zTaAHNbPivjpiYvduEHZ11S
IBkuXiuWalTz736RZxt9fGBqpaREFb95R0Yx4p+G4RVr1usHezWpFvTBrTv0lx7l
KIpTr2C619i47qXuCXyJPDNuMxg5cB848X2EGzFxJ2gwQS9WQ5gVuYGfnTLjI9d6
l4VqUSynHk/OuwMZh5x1+GJTpj8HOR8k3lp3caIxdrfB3PDeYNzMRKNbQGp6rizr
D4Ro99qpCT91QTFoB+ZhfmoBdIY85srMwTAC8UA5mI6wZtjIrzG8YVe9kHk3HTz5
ke2wO1+kVFxAQUUNgaj2Vq9EMttXtU5MsSPIPNcn1Yzh6DGEzEPH+PlhsWccmIB1
P5L117BbYEGrMlA2dr2dkhPxqo9KEUah2WkuaLiHAsMqHFQP6RWtxeB/Xy+r/JiD
eBL4ATHHaguMbg5R48gabyMtsEDDobToCSNyMZ3mY/c9ES3fpLwNCGShrOZcDRuU
z3OlZD21ogUVpan8wDkEiQcCUEhadT1FdcVp9Bsa/aefYLXXrHj2C72RJ+gcJLjt
urRQme065ivK0wGRZVgoXD7sNv5zyOwF5A8wUhLuNyxvmCkGu1Xo9E9JUct5ZX1j
Zc9qhc8qECXHxy8iMezVmItBKDKEKEMIQ+SqbYk+Xt+rdEFLuie3Y3etLkBuIU6r
HWeqImqrRSJZ1gFKnbyQRnzDdtqCWpVxcWkxsExG2YXbdNjpUojuYUvpvOay+M5Z
pVCGve3rc6PbcncRr18yIe2lqtDlYa3KW4/AnJIbOGPFks7CjQpm1rHF471Td8u8
FByrbCnk/bZ1W5ToTwROFdN8j6mkaCxsOXB3lgnA6gZk8IvkCv2VW7wDdY2g64hU
d8ZrCL7+4COGlnUT3iUbSh6s9F5K+3YPLF3hlK/hPS+Wgy04EHmYT36+7TbrTEOx
W2aLiiDi9T2ykJHvFWdrFZRFQfYrLZhtWFUyQs2RNp6/NpL9Co2FirJp31ElhrZ7
g4ebGBRAQ8JLqxDxjQNivqpnxwBKffUvKphz4lGO18GzHXBvkQ4aLQLiGS6kAdw9
Zr2Z32c/e8wBIB8lqh4QY4L4gv0VVggRSo/pTSO5CRIWV4nNz4ihhTkbjj3XZzr+
AAhclt6ACSYhzi5yf0YwwzGrSC6XrV27MdIP5gT9z6e5x+CjFW6rg7EFDjQSoDEt
l9QguIlNd7RGQE2MGg9Jm+PkvNbEvFFW8HVLsPV5vPcrUxVzuL1gEyL/mut2fcYW
ZMKfvtOQqJXjneQ3O6ofE787tXwNUMFSvvgO3x+YTCtomyIzlRlLqEuysEObab4J
jOnnbVMn/KX1Wh/EfuNaa2JRP3dYBCZFr2APMGwcbAOWjBgtQmC4W2+jd4DDcotn
Rd7DuXZ5zVevWsE6jESTPrSpYqddcTGj3wGVDEk3jnRDd5uT3QDCpMXyCZSQv1AC
Ln15Q2ksnGv7Ff4Sppa4PgtuHGrZf/lRetLGoOEb0+Qa7XQThpamBhAcPlFD9cja
A912FsB1JxnWwk/gKVMP6D/2Xa2hlMSnbCjRQ0Gyll1N5xV2ZOeYBHAbuEfi5sYT
UEpdoGjl1EzHfIyP0dmA6ohOFKb8OrOBUXbG1fHOMqEWx6BKaIE6P1ZwJIGr4k4h
h3yzS3Kip2hmMVc56BwhSfMJM2srlaePz8o42TA4cSwQexfpxv0apck+B9ygC6Yh
yY55IGAJXy3bcYTulMBvIFxL5MJNOj/tP2G62Z3LsCtzlcdLAdiKlcuqXCBr8CPQ
WvLRV8TaznmgIc4W/sqbLMkcprJtS9RwA3Zbn/zeCghlYYGGYbfgN7YXun/BrsjG
VcZ3pghPm4HnXWAkS2sOxFvaotviGE/fsohgb9tyD8/COQnTIOmKmPpe9u6Ghap/
mBRovAQYh720IXCOHOkdXUuclu/7QRwBEv/mk2xVeltgOnmQMuICRL0Myym4XWMP
U4j9VEHuFOFr3aXVCboFY9HLodzkM+UKaGB6bxIoOixb+C4EGydDhV3dkv7tdOF7
dOzQrcD81od5lJDg2aIns3nbDPE/n8uYKGrQ6sdlBiUC9lE/Du+JSRwi5C4iJiaI
kFG4I03xWH09y4Ho8WJ6XGOJ1WyRTXtnCVCNOdh60AWFGAzVTLs1cxpKSnRgKZk4
TusWfC8I75mxM8LjBLnrnFhcw+9NUAucvoRnGu7xmEX8YsV3Dq/gYB7VUmqowi3+
+81IgmH5HLvnTkmStyLIMIrzyEB+h3j5tE2u7evw7RGpJjmt7f6kT6f0iwW9v5tw
jsFRy8f5uGrziUA4QMQkn/olG+BsSRxLkL2YMM2FtfA3yVmpA1DyyWWFTG1lRvtw
JBA77n52dkEz3BPo5Sc+DfuRPnwNHKzEd2IFcMGtSAgWnO6/T/V3E806XBupyU3z
vpv0zxvE+3p9LW0J0Z/RnX8EmCQknwivLF0SC6CIE987NQh+S2IufAF6yS2stF8E
TmP4OL5xJZkeTEZKEseE+YkA2B1YHXGfLgDlWgJ2oQXZmC2y08hTyfuDd3zgl2Ez
BckJpVgxLGLgM1aX3MianqWHpPA5zcprzFQwF0mr9aDtzGikeD7lRSNqjboNjwEg
egpXW0Y7rSa/GCWl72cI+nY9GEYpEw4aFVzgqbPUCGNon0dtQFB+PiqaF3dEvnLE
R9qCDkQDnR/kU2dsRB4TOOwsZWRZnt9FCNSqEU3lPruEH1v6am7tmP/kni8a8pqt
vJI9ls4BdrLg1C5e17ty0J+16C7sSuCyMUWtYg1CbpkDoTTf5TH83uxpKDaJTy4o
OeSPnVApZnInWyOlgPpwcEDDHrsUlkPvgFLiKRfTTeBHUptuYtiDxz8MWlGhy076
Dw+OjpxZNC9R53wYe1ct3yRLdvyDhGK6fz6ivMjFy8HyJtWZrY5SWFUPYVH7TXmY
ZG0w3sZCLgHhsVnqDZo/NZBoNvK2h94+RfHuHTdsufmsHWhFp6O0b4DP7mPH8USk
63/P3OLrGuHOJhSlDTQ/s/1Bf6UGQyU20WYHTeIOuXO5zRp0wfjHpM1lNEIEkcOK
gH1Xu4imDaX56S1sVS5zB/NPLSBQ5nUMkIqMvEZKYS9qZu1fDD/R3sn0DXtq6YLQ
XScmIfFXIa6dXRswXBmjzg3M82d4gRCMoXtHlmcsZznYoAlyVDzeClnOyaQQPJqZ
TBadyEVimQhtAws/i1WFapju04H2VmykDlS82s6Ivnz+Bxt0ejeLumCZm3Q80EZT
l/lDlu0EKYWWivWLOBLHLmQ/AP0+5hGNEQC58J32YJtsdQzs6TlPaKAFMbR04LQE
ZgpFxZ1mT8V+iWdhNhSTRDQqFjei9qHDKNDorERlnDbO0EZP+fQS0b7akMYhd++Y
zqz8NrnY6+yt6D/9UDWPgSKblfPao6uRep1G4q/K49m7lfgiX4ERtTBhm5vX3ZHX
9NrarzLGYkE+P73vGilki7pBvXAX3VzSm6nCi9YKnbh9qzqLDqA3+RxNvS19uMwB
WvQ3eP25McLBAzElRoB4LGYDkb9HiYZoXIkCbCSLnNN8gEhW2dufB1rD1Hvp/n1b
OVksmlRmDW27Wlocv7YN0OHd8yuSW4KOvwVYMty+4bhdGd0xT5gKoJ1Hf84w/zsx
/4vU+VgfZKdS1ZtlLF+Qu1zi5fTYyszht88WMnH7MR9P4sq3RD8KkwAYKa3yZJEJ
cUnqrINjf2ZqAUMDq+L5eAF408vzn3AojpXyYCRW6zYPmGrZbObNygbHxSE9RbHW
JgpmFAnzMbb4CEp775ezCQUDrWgS2VDS5veOaoM2WfgQOp5/PLJIjUDb0TwzBGzP
0CCKQA/PIt91htul7K94CJq5CvIJ49aTdXLtLmtLwKEyvADkZMy+Pjg3m0OKZBXY
B8BfVMGcAhPgUF/PvDOv7g+r7MEc46WtkRB/9DxhnxTvBODXLxjRiPmBdozRgZuZ
F6mP29zJPQ+Us+CaC+3oHWgng1E96dOlyg+JISo1phcf+8L2f4V9sNubC3NVb8mH
o8canB5ozP3uS+NiGw9rL3BPqaj0MNwHz8azUueJ7d+y2cIrWiZeQ8obkP1oYns1
hlJvLVn4gXjTQD0G38kb7fbLYP4oMuk11YmDzaK/n1jcSt/LDgr9JKERXdOmpQU3
b2COdVOtTeR+sl3q5FXyf+nZNuuA+N1+AGkWI6trzfh93QkMuDuoLUsBeVPTUsiu
Q1D/DnGZrqjACtJJlr/fiQtttj3IndJaSQHn5tsaB2JNl8Xll4HCN5SnAjVXqyY4
TxFlvAaEyx06Uho3cCGp4UfAQbKLYV6Oud3b4HXYq2202VMAkF+EEAe8oPsFoLLQ
qsa2GOl9itGGClDfy3gg2C4nYil68F096U9lCpWYls/cNH9YsqR6Ic+m3GpaTy5v
v2gvIxZbC1IHbe673FT4NjhcwHtZSTA61gSF+NW0nZLVRTudqs+g6NnvOZA81qi4
gjkTmP/vVMXHHkBnk2fvOmj94vNOG3BEfzSUKbaY1lZ3RVJGx/j7kvCXRbRVP0A7
bkWX5ahwNDXEkaHMy8uUCc4vH1t5ETkt8AjlzLury9PrF2il9VdBI32JOfTfp61k
P+wLQCaaaIAwLJX4wzeOeeL1nTVOoZARt5Sncm/weo2fCPtdKjt1cpD/0aviZOgU
HG5nbMMkZNXkMPHmNeVb/xvwT3NnRYYT+R5FHYCyJby7say0uBmBcQTHkEj110RR
/vui75R2UDFlvsf6nq/CjC+gtF4pPzyHmuXwQnNdOg6DWOJl01iq25xy5osNFeNj
g2odA+mZaOWkGhTk8BdQqcI4RnUAJjJRjhp932eHxKoHqqh7OMyg3kfI3jo0cW/8
4mILCPT50zVbS3E1+KFJuR+RRdY7s2K3ObG9pIk9Q3uqtE7KxAi2BVi7N/53acho
2lxFiqCgyLjOqSHB9BDYyq3veHIPTIWq6p03oecWVOIOCosHvFC//3eFoheBW/Js
TlQ1kypQfdk9o1EjlbCN3RqzTjDyQZ33ZxmDsQuxCI96WV24hjECHk/vaglQFeP2
39SXLDyEjUkOGgmUyWdHjqMr+619RL2lYP9d1USAn+z4IVTfQBlZkuMebqm4sms3
sokH7aYRxVE++bC3qZeDOEbh/iYMpXPWfkB/VZ6Dq7GvbAP7V4n9i2scesHFhEiI
D55H42ZGNyf+D7tsROs+k7tP5rQsCq+badUsm7e5l0VOwl5xNPHxpyITH07KZzBf
OyTnmSm685CvxaMN2+8TST1HOLeZIfbHQxEPsaF1hMoQHq/XXZbDh4nestFQBo0q
w4lNyEkieg/TXh9eMbkUrVX2tFfVUKlGE6etnH4z70aAgGf0ckHw+/QYAHyRSuFL
UVrQ4Av6WrsVyQlLjKxzv/Ke9tABRXfk22jXD5Vq0hRNyyhzcNObfS6uayUwdozO
ToNN28Ymc/cu7UGtOwLMKKIRX4mvrkrPZguvg0+Fahz+SgwqMprXZsDSyqmOfoDl
oRHNrqHNDfw97fbAYBtmZmVqB5QSuc8QyR3SXez23j9CeA0WWdbzE5M/H+JqhFd2
`protect END_PROTECTED
