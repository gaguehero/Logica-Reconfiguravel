`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WVvUyuV85qW2YXVVYV+NbgxdW2si1mETPwRY2DxXV+jA2XwlghIXAbtVaw43Mx0o
R9WzH1yZI5PYC1BMudBwaDnaV4uLtPPTIMRq8zLhiPbqRsG5BJFRz9/j1tzvpU6U
t4gpPwil/mPWrGBqKUp8s0m/R9C4XqX8MVVyJPO188bOdWdgcHucm+dFXg4IypxP
7knLBFRG1mKnneFAlVTbjpjDazvMzUM2LShybzO8vvMl9W31PKWgp4spKzZ/taGL
Lt2uVNmXCTr+NlpZT713x95GtlZ2n79saw6ne2L+I6OUghDzpSZG0BcaYtsej8v6
+FLIe5gOYs7FOhBppRLd9MY/0B73eULmQ1JrZOFj7xDGCknmExgQsTw3hLBngzuT
ejT/Ok549Br1E3zE14sqpHPvoVA+2OCQmSukG0dYc9Vt9Q1qFEDCaxUwzMGKyiRE
BwFiJHaSX0W+DhWb5uEReDmr9rcnw4qUZD2i9YINRz119e1FgVNRK1I9lJZ1XKVa
PLh5/u4nAnSQ/xXsLhRmqE6FRAzvpebvM8lPiUnTAnrzjal9ceB/CNxeMQA8Rygj
yzPcCCrN5JeZkLAdDDyqlXnjWW76eU1pXHMfYzt72/OyF0ImxgaLk3tvh3viOHbj
XF3BIZOrtno5nQDuKXP96QqSlOxJmpn8zYc7fdXf1XlREwCDlggl/EszlpBlb2V+
nymcVsJaXij1SC1FgPlkE2djPXk8vU780ChxuQpEgIeOuWHaC259IDGdVPqLNsi3
z6IPoQyMr3YYICz/dPmudr4Ozo230BrNY1UMrWFYdVGhPxPoghFiOxZdQiByz3EU
N3fR26t/jVpMggk/eWJPvkTP0vECwt/+IsqOpNAXeaenLvVxSBkEeqZw1um0JsOz
rJIxmYcTZKSUrsFdjrDyfaxRQUteTrbGpjrfx6n4Fnnra6F8QSMiqX6vt1EHVBvn
AHfayE0dODVY6BpriQvCZgDEVvB5b8kR8TGQZ+pbso4nXo545KJh5LzXpkN3hgJE
PPNo6sFkVxtHg3EA3lQL7LkXtB7VPBqtqZO2A+M2O3rnhgVSoVpOV9QhRGFTmmUl
WwMVzNzPLkptAQ+piIGJsfCixNqRTTTVK9X2QG21m5mo442gjgqOpS8yykwcMTjs
LnK/XPjgDvGqWdF0j5c+aind5Uvb3Qspwbr7EnPO53wzMUBST9obg42MuRz/gt6v
OicTc2+4Im86sZNhZ29s/2ZZkkfjLTJCfny0vvPsiF2BNJ4Y3BRDJkoVY4cNrPfB
oXt2Q9hfzp/rCljcW32FdrdTcNUDuzm+yoE3wPK65ov9Ot5fNfFTyTbg+BXwn7Re
DC2WdnyFjDwjZQCj+9QEoxE2/61IT7f62+5HyYsK25T1dEjCpMsOxB+UF0h8dPsc
ksK1VMB/cO8MzRUwqDtNm9JLT0C0fndYA7JlmVNhbRui+T9a2SKTVYSeIKpNjh2o
H7aWpo0h/O/t61YYxMx9aiaoWjFja1JtbxDq6tXMAIoAs+Z5kOzFy7KGw0nOoTcF
wucXHkZlArSYM8Owa+wc02G3IqtDK379oaK4iiYwh4FbkzNUHUYPsHH6atnSEHO4
62VvzSx8TiGUgHhLSfi2IuOyTQSGnRDHE0ScR1AeBjsjT8L1Hh9H9WyLy4O7ACG8
wuyhyy5lAXde3KozevbErIVlDkYUzqPDNWleyk2ZCLDqv7Llfpf+uVxwv7F8U24F
JRfuA6Kw6U5Gz3pByI//HrFeq7+ixlikBjsinMdn+fKtNOO2A773EvgyCuhF+8Ku
u2keFUq072JnCFoNDuav1pNSCqRtvudR9Kx/UwI0dRrKYnXVlibZToptPC+88/OC
miAoR+VLiy1NngwjiaCU6IRG2eTakTP840tZ4m0BBV0gU1uhZrY8LzZafpQiIfE/
xNJY4Fdih4ga5LC9J6P1HpD4lqr92lXI/ij2TNuP4R7uM0jHwfjhqofIFqgVWQLW
KwodHVTwu1y+MlWFO1hF3h3R0nW5VInzxLOKRH3sAXfPodi81ftFx8k1GTzLFhH7
Co/PhQUlFlLcc5pkOhplBzaENu+Cnq5TKo6KqN0MgAAMWOMQzTgA14yMKz1SqRwJ
tr92QOvcNaMppeDZ1Qrh5TxA/PfxGmZJr6EUNtxchqzo6BJC6lYMNILkyJ0jSzex
muRU/6Y3gjZvL7BtaWgaJXe/iza0fiZv84iKNzvFNrNP1ANnn42/TG/RS8QF5MrE
hZ1NVc2zJKozLNM44yv9TQyfdJlDqFaB04K7hIKam0oLeSdxttZR2aanBR5EaFIw
84DwJpAU6pqYwvXjEtRo7SSMRGNfTjV8Q/uH52uZFlcbCSOEC7bh8hWmeYdqxNDb
bs3NdgOruAzBUryxBIYeq5q4mD4CXOwdPtsrDaiyhDeOS2oT//SmmEy3gPYgvtD9
EVqmxejGhQ/9fmV73ozRKSZMEvLLn9L0ZVQ64JFg2eTG2fMY5l188Jbg8wh532jn
kZAdIQ5tCiDZl0fERAw6ZDMnANQizhc0poQnTrsR9IiCrUrcVm9wo5arXXx3TNRa
/+S7sGIs/xG06EWSgYTGhmSYdZyK1zxcLfybOmHnafkz0p8sQ4GuBFA2nzVPP8E4
368Exgv7Bpbdc4VcuoI4bmTIsVChW4e9BZkG2rrCupEh6potIA3RYeHzElxsWtsv
G3kPi3nvLdryLoLAALiS1l6Pb18efOW7U1Lm7748OkmODfNJ6uakrfyQb0/ek3o6
eBCLSySSg85EuSwI3lLQx+209csoNUMGktcVtYTE1bx1A4hKlKGeWhug0sYJh/Rz
3Qmn2qyBFEMxr69Sh0FjdbuYZGa3rxqE1WryheluPWKSBfV0/Mt4WijUm2aExCN6
LVstKp7JTeeEHOYO6hR8JTLLAbk/Zs2ctOY34hY0SNMPqKIyPHgXhQxE6nban6sw
T9HWfgaiEPn0XAPj6He5Ocnjhi428x4MtMSLABd+22vXfTzNHFKm2SfRX2saBjzD
nzgPWWEjkW1c9OMZ8y64M8/cy+8e6pzUHMSXIcV3gQrjzx5eX4yqPfnC+bwQhtxW
mWb32VRDyNbs2QGTWL0bH0v1lNkcbIYpdh45hF/KAJTlhcjlmXC07knC83KF2B3L
et9pwC+goIeEEHYq620qCbx8lytz66vUgAmrBFssNltDQjDZ36x5bxXdEn6p0KL2
ei3QaVZR8/QyYaYuBBuPvxCpvhDHF+XELHmC2d2poCEr7TK0JpA78sHAv9HtZtc5
C5NdyCOuiTJCklYyOHgKPQHINZQq4e8Id1QruWAn+SptBNpa6AqU5jal92kxRPLc
MWSEvb1qBljvj5XXn9XxFQFuqG1yC3JkKwwf3KJoJxH3WarOLg3GMOmHgZs+2vGy
HdFUYu2dncCS3m57hpx74UXQeKu4CnyrNQn7SIadVSfuhqe9o2XOQd0dpBrXCQV3
lGaRZIifJH6rysW7uNKXBKB2kcEtzWqXl8lAImDIlc7xoiLH2uMrtwxwAY0/M3FZ
5KFHwFsdI2bkorDv4crZOMcmpyv7qs+0m8FGvQTrQL4CA7OzOWaFVwq9sUUUjnfD
75uTfHxoBb5kkOhM1zBjhz9qcCicVEB1pehoptYVzx7jjfAuAlqDRNfEeDtppOwH
zy/QQqvAroHlEKtR/GmQ1W2QS7p1VIUkRRJCrBAwYWBTWAs6JQ14D9U07dXbRf3o
6FNUMUEtuYIPrQTuiexLn6LWPC0sP2tvzOlHuLcfR4sWscYLWIjpM55Y7pJr/AJj
nNEUG3KjvuhSJwCTtiMXgQ/YkzjYVUN4itKUR/mXH2uPpGu+AyGicN1bjghSB9vZ
sgr2Qmo6fvdHeVLK77PJ5UFe/HAwocPwj45/AnRo4w3JKzVaRe0iYXpniyopyiQO
qTSvHHn6/g7D4AjakEria9O48EunpAcjkgwmQZJD6VYjyRi0u/kr9uEhOgDla2OD
9/3G3Mssb2VYkqT2rMtIl/EotySLvgu1fH8Y8q6e/s2sjHmRkZ16hrJ4T3FW0HEv
ZkAEPg69nD+qt/46tmX5GsTwOtvNLfwd45R50cfcdX7RndXTNYpQsaP0Wa2M/d6p
QqZUTTd0SVmnqVqJ389+577iuoj2u1QNhayHTao1AVf20+1hF5Jlt31S5gzQxU3F
Q34ur8PAMi3Mbtp7b8FN55E7lUfxVzlOYLA3jEXWAZoGXsa1kL5uNTvO8TqgUf7k
nbD3YbXKf3/GY4qwNBSiLtO4WTxottb25nqXyjp5I8ko6q6zNufiQFyPsCAY5P7L
J2b93+HvP5AECrufyoeCyuKgrlguUnR+qtRvB+acfppoxyEhLQwTSePhbvQbZokZ
Iqr5Dx+v5/JFC/Uza75zjtE3HiZZW9SAMbgGAl9Mz5wInb/ZUa0uMJ5Brz9Qkl0M
j8BguqkTbAHH56W7oa1ZtO99MEloQEDgZ4K1+82ZMWhZzod60fiI0rVBjRdE/RGu
wx56eFGGJXe1DowWY8SWEk6JWu9eQTlrky3rW1J+ABZPYWBpCDByJvYm16hkVGXt
ACOuq+CYIHXnIxMVWPJVsPtQxi054QKtDBVrB2yAHUR39x1R2RdtWAmfBGzlG8j0
IIg5JDafJcyQgRoGG5S8w1CjumoC1+VTKWBBRvn6B1tv/YiZn8+G8dR/UUu94p45
4VfjxzL1xKgdcEw6vr34zL1YT7TKliF69Th1fnkVa0zfNr+ENFKMpA8oOel48s6B
vL6LGwreZTXeuY+UlakZoZcMC0ePPs65JEboo7lLqMKezwswR6o6cY2edwtVLOu5
xeq/T7x7DFRT+J+h7zl21NFrd6QOLQkqGvypQ2OH9g49KR0VUYKqOHBpto9N+Hok
tCcxBAQCAULBTtQj7WMcp8k9zdvrwfTwLf4isqPdAwmyaH6yIRMJU+2rfDhVqAHe
HU5R68eYK80T36pBDY9Bhju3HUxCpL5YOFASZnrOGj3RBuPJ2ErWj4eH+gkGda2C
dn1DDLGcSG4UOQxfC47CuLkZMS6QgEad3upmx27U2JZxS6KCg07ErPZmSgjhUh5M
ghN8PhiVVt2/N5lc5j7OaAbrUcqe2hcmXR8JdHDA/MoVjYHo7jThzQhVsmlRY7Mk
X4E6yj4cbzDNC/LK1Aw7bjZdn2SitO/bE3cIvkKVP/je8zOD0EIlj8xvQQgJSQtq
5TrAmelODpxkFJSjXEfxR9lABMlEJWtIE30VQ2Eex5FcW9w3qZgJPrXIlBI/7inu
THJh0FqYKmfdDMq8N7kxIXif21fXRmcJ6ofX4N1Y4FuJjhaX8DuDxGkBp33GCpfK
ShTF4zURx63cOithPBGO0mhCHWpOHMUNTXYZDu7/0s7x50+12LVPml4O6gRcAfHl
uhbJz3awHLXML9waZKGqNZAiYmCFH37Qrp20Q6dd1LFuYbjKNcms+tp6PrnhEOWR
fHmnx6oUF2t+KDt4BLMCF+wGRKLfx51owaYwbevxo5M+NQonoxgmerogPCMykONn
x1H4K8lYIeO/bnD0zC7mhwemqYf2fisPA8aPr+coa+ihp7cYE8IO7S4EN6Zfd1zn
4B5GU83FWoC1Gld9uTvcWijkeTmVyW6We6jjTMRbNu52gKt7FDpvNyhKo9lNLqZA
dWz0o9sOgoeyChI/oZxGBZA8p7uoD/esGkghkPJS7XQYY1ILnMIHLb7fWFNvo/Tj
Az+wVo1r/u3zvJNVYXy2IE4fj/fWMp9kajS5FyuGH/VWpC4fzDSJ60ayFfzwkVCc
Y2IpfBrQFvHPjgpcLbFircGaIPzQeo6j4iJ/vTd/rqhNrdPHOS3vVKuNlKRQukkK
5G5UdSWe9fGhqXRhU9vPA6x+/neiTsScLj4UJDErljJM6rp3V3fODm7a+JGudCYL
R5klRu/LS/A6cbpPf53j+DJ4cFQkEiHaAvp1mD9SQF5cyl99flXJIH79r92tIjnv
VUAwM9gwWldZRiLps5dS0alOEbH3bnmtNApZj/gx6/C3bO1B/7mj7hWcevcREcle
BtlnUpWLS+4we2KubMlpq8XNP65g8gKLIss3J9xEGfStyLtVrTwB/ezHAmiBl3Rt
CfP2Wu9hTyEYRELBp5P+Bb+XcnajRBpWxrIxMMg3jFk4bHL+woV5Xt2I7aahIw2R
m+Tvgn2EJnxdlELPgJWNeiNkxhvTTlO/6iwrPUoN9HiGinxXvq691J3wymYP1ENa
AV14QCTE06aHVb1YVvwUDmxxCZzRGru7nNrqv+UqfVtupdQrDSxKX/fRCel/CTm9
+hloss2n/XKzIkGCP7O1btvYY+qvJnzSzMqyVE7Zd5+hRx/CZfnD96dTSZ63Tar6
EP2AagBzRdJbNOGu13kH6sUIuw6K8kNRPIYy/LDuJ4ZIQAlYp7Fs21SP5EOTHA5/
GluN4NGPhoUks7vrIVXRlVaetPbiR0ZWcSD3oSKhHPUw294OT7ijWW9YaoXULLze
3q5/a6ivPqGfKx87TZpYSEJ50zmdcuO3IQTbtme9E4YKVVoRBuSDxW9jQYgFdPQe
Bjbuv1B+QBHRdfa1rKjcczR1Ih15rh4GnMsXhAHmzB+lssHZ/KJ8RR9mw6nRNc/0
XaSlN53F6IyjYyd9YwdNohyHf6ADkeYE9p1tnMm2me2KrK5mYSvWlD4bUbhCJwVq
rCv9WjsuoHDD23FQkEr77LI62fTgKAtlml5ZutIf9EM=
`protect END_PROTECTED
