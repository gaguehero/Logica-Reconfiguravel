`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0scsh41sg63fXVyDHl4V+cW9TS5gmUFYRvq7Xpa/ocDuHdk25Ih2Dko5qdRt4hF
/JaKzGXWEC+Or6wtGG5qVXSMnzVLNuKaRBqqUNr4zoL/lFK3Li5dkgpTn3iVodHo
3/J8HO4DUY/0vqqCd2BZk6K/aVn+3XzJhW6FDolS3AdIQ9MKPJNaK3MLDzmQdfIB
yX/4R3oH6Q63M3i+Uta/V0e6jg9JHvYl6lct0D16WWPqLNwwJe2usKUaWpNj9u3P
bOkN7lI16EGxnzONO3D5eVFplYzGsOPvb9aUJhjL2a8Od+tMUNNWgFjiUkHRUVqv
OKtF94BlmZqAzjgWyHHp50mvrqBxbO4M5k3fhyYQOa2UF53QLsNXJ4QOs6UnNVmO
kHzD/NZU1Qgjabcxbj2CmY+3ACsNmgtxbwW67Raqhk1QF2KnYSJCfJ9TcuODDzBn
fFwhaVm2JnckMvNCBpRx3udcoPWjuUhOgh34iEQsF/ko6rVEDPAEINxX2GBB+dCp
JzGGv/1S1MtLHsVFqxAPYdvy8sxc7XcpZbBAt2eH0c2BNGDcq2yt2Pdj2RTdKNlI
HpmyYg7N0YTWu40KvmWXb7yp9BMkUnQwSe9o8+RtP94=
`protect END_PROTECTED
