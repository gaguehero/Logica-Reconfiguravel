library verilog;
use verilog.vl_types.all;
entity cont4_vlg_vec_tst is
end cont4_vlg_vec_tst;
