`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+wVAxJ2VtCKvE67XINqCpCD5WxtZkqga9Kxw/d8PlIbbc+dFhsJ6IB/T3eJkg5x
1lh0KmwIMUZzDL5rvm16NLi+RTvUriPWr64DT9GAP9Mg8AAq10agqflezljnP/8l
QbSBKVbgAFIegED0QJJdd3SLW5CUJM2qTfBRNaZfxin6Nk/IalQZgDE2mICRsuvU
OSFUr2WwB0kft3GN7CVIrPhxlv0lcYi1oI2wG46Y7SPmIZyLy9VvutRhC17putqR
S3eMJY6WfDYcPO/EhgCD9L7cM50Hc0zGLUNYvTULNv/rj6AnPFl+aqCgFMooAMIn
FCs/3bfqsu7ReMs0tDiRSXwRRJlofKHC4hoGrNJ5tJEFLahtERVCbFhH7Qy27ykn
m8+XvYtGiQyVRCkajjwZvTuD1V+thmMjPP7A2psQWVkh0ZGdV/5S8DYDAgw87AvZ
TOpI7ec8I20E/trOjrsDR3Au71/JxEWW9wLbBalUmRKVLZIYPLNh1y3I9i8au5z1
OemjwQ1jp2acyRdtHsvgRTQD2pxH1xXMWfbhOVpPcSXe6bkzLEascZXT2FGeirWk
m6yO/IHmMu4K8EVisRMiNtXAL4zNAIiYDyzkD2v2uLhIPWRLXsTkP8B9A1VKlxPR
P8zr2iDd4e2eiPt6MX0ooLogxeuKI5qUE4xRREwvKusEk56C9Bn7zuV/HeM7CvSm
ML2SVQCPluToj8DzJoqzyYCQvd5wOQtVzp/DRUMdW4aoSuYVUjsQ5MuC4gSaItVd
g3WrK/HTMCYr2vwqzKW9vXIOsVrGOpDMW8E/3qAbmIFZCMIfhye03+cU9m39ZFtF
ST2B/IBUfQ3b+6JuHWxDaeFyo8aZszWWQdfVSQsXLoWQttbLWB1AVjMJHSDwnGI6
eh2N1aqQq0PY379uvTR96HBijySk2rOQwgWKtVLW6081YOMCftIQzHA1guXOHHBb
IjwAW8ICF7gnwxWmn5Yw0ycgiO+DpTvUjXQCxpU/6+vf+GLSlb112pT4ia2m+jeb
WMLQ520NGkg/X05zfogT/ikVXYa9CAu4icOdpluY86mJwaq8ZMLONXZ6uWUNklUm
Pziyp7UPqj8oSnu8Wmcvb/kgU7/HkZZhdDvEqiYbVVdHI3qe7pkjwbMVDm2icuy5
s3PWcyFFPrJ4z1n4XLpPaadUuaLrUKAltirOQxyT+6+4JQc6yXwGBvo/dik1FmND
M1czESicClkhO56YPb0bvYz/LYhUu3pM2CR9nB3jPR2ju8Bm9TxH74fqO9OutJL0
w3PopDXTFlW7QtnHAK0IE+xBNEno9cMjDtv6euuADBSOquZdcVpWkRl7DlC8Xssy
C0jsAKOZvGCoN450hlwq2Rej+eCgPlThs5e4gBXxCS1vWJgtOaeXMTf9zKq1SG8c
7s2dn2g6BRpldY7jrIF4zE8+vOSbhYfx1NqCfiqNUNQWOPmgzcilJ9peOHJBAeUH
y5VAIxdG0pEdjnOlRFlatFVe3WAb3DeedCQuw5M1w5wecEK9eA7xA0Y0qUQ6+gzQ
k5uGN6iL737a+Fpi8TL2fBETxY7SDoQN5x2NpPm5D5Qy4X82HqE4P0cyAnYgqgrK
CgMvIqt+WYVeHRbksFhEgXdnuOFPq4F9ILLggxXsH04CsYgr4y2OMBKlNdQL6RLF
WwkeANSzICbLSdkzO+dX1ynCHf8iir8QrHhy5syGuieoD9VT/NZlSOi0vv2Y4FZ7
+GJsCtCVrf5eGEQFmsxHk/r5ZMp/RB6r3cNErIoxhf8d7PumIXWFZIB9ajgLI827
VLWUCDP4ZPSjueSgzPadUfEi7V2uqMCyJWdZlkMGDwb4/+RcWyS0HiPnDTHlvqfi
z1MgC9H+FzWV9XNtNyVLIcr4PdjaTTz0LilzscIked+SqM1hFLlDPnALRqEY3Bvm
zVT/CFgxMEBu3PodRT9y8hn4XoGnej9xyCy5oRhnUkQo/YUueL+JxuOy5DqNsRxq
WdpwfmP2hBvQxdM2REhx3n7hBwSW6+6sYCCouCnJDgr0asVykHPL74wbzQfjOGyE
sej53Dl/p1gKw+pc+BAz6Q==
`protect END_PROTECTED
