`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yb2O92UtmiBnd4s8pDUN5CASmrJ3vh1I/DpYjtuYkj+0vCiZADVTv6VaArfqMqAk
mJn1njBQH7yxb1iC0ABwHbINSNgl7H1/AiQI6OoPqW3DzdI82thWwg8qeAhf9/XM
REiEqy4+Fu0zaQ91HFqA3AjI12OFwU1zPCR+FWGIPhrYlywvZVNAXYO7ieRCY18p
HPd5116UD8bamHtXYjW7EFmqkpBXuRxaOpaDzzMqpGUg8rLm0sV5DFMy0tAMhTGw
9gPGeaxls5pzEhzwgeddT+BGU5rR3t3f0d15sWU38QzYCtTjRNOLYl6fwmVm4fxj
oxmhvlXvFF/v6R4arWu7OMJbkWR50pEWFiqICJvYecCw5azgsGLT+moLSHbmB2Jc
aUyxFlDdGTwctWvH6kRR6C80hLDmrk4FD5EfxCBlVjYmznzgRQ4Ir4lhHyJVy9vK
5XgJoLGx21RNXOOVWJwiLDZ+nQj8cf7ZB9wVvEHUyqdBo3E8nSkWjBbXWHaD84EV
RK/+4vqNYQ5BZ7RwgcqBiz6MkblGIsOu2MvcU6R6U0q1SV/2WX+2X1fO+UMMGljV
ML0eQtrfL2HQsVCziJFFfUC8WlO/xkaMPSOkRnmw2Fp8bxoddg0sBKlU7tmLUREc
+yB3QFcIwizDmctioS0AHlzvj0hMs7EVlbhEHvafWB+ViDJJU1ABb1VBQmh1I96K
OViKYNb9Aun5dNoc8tw3f73wlkoG9dckD/VUNhAuU05BTUrmbP/ovNVHX3agdXzm
/S4DqnVeZ6Jm6+OI6P9MG9Eb2zTm5ouKR67KUp8UCbTSsfEUgkPZeWdMchgLH/Sy
9zI16x77nKoUUhk+Zi04ZI/hKng9O5xWmAv74a2gyBTsn4vxx/ptp/MHfbI9FXQV
sefewx0v/SnJ9y09OEJ8tZYzBPWNWyZcWjyvROVLCl65Nwq+h+7b1U0be0T91r5b
EJgsVEtiP4PhATrQ6waRYekfFQoJqonYpNst5/ANoEnAJTkqzkZLpZ/VeKV7hnQ/
UJc+Mju0dmwLVKUQ2yfCZn6Gq9/rr7U3yjS9Uus5bx2rVZ3xHLAbKt4d925EW6J4
nt9jW7pm7D/81wBpMm1OdKdnSZV71K2yLxJDZPLh/PHKmLiX1Qjqa4AtW/oljZR0
FqLjjLPGVTH/WVqZUHW95+S4HX8jUiN3ezshSTOoAlf87BydvjavUkom+ip5Uu/y
CKIhqjehXo8EBdj3VgH9kBjQNXwAgkCr5AI7afOKW5/6VvTy7sjX/RZs6S6t2PXv
PmBsE+ceQbz1t6HXnhEqjaKX1WcJWgzwvrl+IyiiEuaMspOHSiy6K3Ocki0IPs0+
C3+BAP4Zc/RgU0bKIzNiIIvY9bUNI2QsVogA+k6mWsCKuL21M1bCzPt1PZyROYOn
L9yCIF650hXD6rZOhL6svWsMt7wl1qKNcWOTe1wwd/XdijTlhJ1GEdkIE8vQ0Lja
MYXQfeRI/q4+dnnLnxqNSgwA6lmuba7+jCy/hgYn6PV3vd/qwwZnYki863qycFaZ
1rXgGLTnO5tm6SgmzqAHcK4Y0FEWrHMOlgnwxG1gxNSjal0Lt9jcNojfDcvcjhSZ
tvbQuAaeWo9KdNRQEypQ5+EFfXwofKBnhDR4JUA++E7tXrj0Y03U9ZgwbVovfvwS
KOVnb1vVXUoMGP8Ox2M1Mn/oWgqc72G4MHB+ZaHytsyYd/PRLJYzsmXcYkcS0RSN
AUPkrzyYMFO114ULpzOyAoIMRvw1c5SEVW3yxGCssGtGLhc7pVljNmglf7+9Jb5f
EK4Y/ayb+OqhN0OnsN3ywz+c/RiZrNPHLaLObXAzXg/nv7SDWhNDdOAdBcWA+Mc2
cB9qpxe04E02k6SQ8hWjEBTGkPFmYyQqeZUXs45pNl49b6a3VL5fYdp+sPM4ATfN
8MQnmvGSxiKI2WHhk+C+DRYu6D8n0WH6Bx1EQ5uC+IMOMzUqdq7Vl0QdlSHQP6rP
tBzoToRdiWsguCquGlGRLKFw5zqHcAdHR+NK45SExk7Oeh7M+twvdU84LofRYv0+
`protect END_PROTECTED
