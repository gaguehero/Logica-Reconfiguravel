`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIAC+6iuxElL+52rbi+gQF9RlwgN2VWIStWH5Y04QsrMIQNt6kOlguEA82qNBSHY
i457z6qVdZmYt4jFCXGHrNkQxUa+ZYtlGwySL7ZalGu2Vzv44JHx1iZflMczB9pC
/VlTwUd1hMN2DaHbqXGmPCwLzEE/b2LuarRIi0jIlVvG5aRCbHtngI7Sz3J6i2k1
LR85HuTE/hysLi56E71AKXEiR3blojSHRYKoxYNOLahZTijjcZPTvJcEkIwsj2d7
psCL8FR6/VBs2UN92BDrjktvMAoqhbucuaSj7vIicuR0x0vp7aDzHuHsHVs+Q04h
exE6RB7j5IyN5PeZuRW6V+1IlCtlbT18AUIQLo+Z+u5SZeVCjvxq/pAe5PPoDvIx
IcyJaFxZgF35nhqv9uvlfKFCKYLZW03lm4DYt+VI+5LiwG8U9Gavg0/qpulJEID3
I4egt+49YUnfBQ7Z8WL07dw1bbTlmKWTIKlP2jfsKUC2EMci1iqGero9rXdYfqRb
tlOQko8jkuu4X31K7DvEbGgMWP7wj1Y5zR6qzGyJ3v/zQpVmReJeva48I3wt/766
2TZhVWnsRkeni4pjd6hzG7UcZz5OI27ZxWk0Whiw47axOCLg9C0BRNCv8v7MAY4G
32m7NKMJIcHMezzaO4cz64ZmBUplv68sfBoDCAWcwr3yoq9+cs+0dzvcxTPc+egc
rX67h+r5P7iD64OTKbq2LSAO/IJ0xLUoLF9HDfcB1Jjm8A/QiQZpLxBiiABmpHzX
R7UD7ZWTn12wJwS4UqO8nwfst9eb2L4zWK4fleciJ4kzoF/wnErNr9LIdxI5ALMj
vaA4qLVETgOtLgiEr9TY6OC+j059OmD+UNlZgd6ktmfY9hlaNhmb9umHP8ZCAv3Y
hUk4ZxM8zQju+8JXhmq4ITlwZxbPRB+oHQaI+mF2hv7EoIDVDSobJcz88EFCdgru
5iK/30WRq1rc6aOa/WYFkW2Zg9TqyjtaiwY3A2uAlX9FvFtCSk2bh3QQDliYNQcO
c10aW0fQKGCZBzWXPqpmzOH9HP32h2HPhBCBPzb6WnwIXOeGYXC/h9zjNraccqhk
TQGwoMsYhbjSrChvmMUPSJnfaZ+1hnY5b6GKI9Lxi5csPVo0/LZXZebDgTZxPDgZ
l9JtsrY02gQTupFubYRqRtakB94Y+dQzcry76kWa4V9x2ci2fv6J8WefuSZmiId7
/QW/MS6xI96UpeUsF1kGr4ym8YbVLl4mzc6oDYpJ39sztu3GTvysf67BXjjtEeJA
QyjgoAoHqkQ4BkP23QPcqwvobJG9kpwezCP3jqLE8kzcb0evxy68Ajyoq1ex5NI9
eHYaJzfHDsIWgnsNfQd4hpStXE6vTb5BMWbeFHwir+2JXCHwrZOQ8JpKTtJWMYfv
BFsb29Ez1jRAR3DHrqM/zeysHfgP6TaC9eT8gW+EKInIzDJE+WfHIuZL6TM0fc7F
54zY6yp1w4Epf+/lfyHiRdvi2F+4RU1ITbWc2nLZ3iz6axVwO3iGHop+ThYreBGI
Rt96C/TNXNpq/GiMuqXmv8d+OyoPAo5I2NBPdMhUtQUZ8MH39VEK1HbpdlLNLmj7
71L6zp92gZc9btTG8Rx6luijye6s7CphMNHB5wHvYxV0KPsua+UunkTIcvFrM7zt
e0MiGrbIYg5GH1DyuM/oWqbDFwDYbUEmWEQRYa8euobabgpTwlGBUpJgeFQ7vKoJ
l1Q/JZRHIyubp4jQrph42DXtia7rXjcx3c3WFPSyjkghl4Gyir5Xp66+625+yWKE
RyysrU37cu0gWdip6fkF3nHoAQ08wcywfZAqTeJmz4ue9XoJj4+2pt4+TDAA4sTK
SNRW5MIbScPQPBsj+/w8ioSsWOyrL89lC7ImCgHSA6GxW/bCLLqleK0nvpaL9CI/
6P9MyTIwqOsto/DsUSlX3HV0hh4Sm2LFW3r6OvyusVZvKurvYSEDGEtBjQrhAXla
qAwSSXTTnUvpFJwIf/e27qzdGfOW0OIuJaSM97qZ9I5JAughf1iAiZtHx/h3fWZ5
kBY+cU5JGKnKI3Jnff0YiQUOBakdtDRwGlDmX3AA4IR9aq2zYyrAdFc64MWofDLg
46R092myi57WgsscOBhrtdj/Sb342DagBb6YaZai5DhDLL5wpJcQRXrl0fXFBjKG
ijZz/YBwXpOVpgZ/B6k5uqJbKBalJ862xZGbqj+plmxl0aE1Vh7ZD4BZURSnTnBb
wmHihhDV/eR9m5VlfxKAoIeg2udUZ4a1SU2xd+zxsNx6WweHvHh6ODD46r7gSHYs
4ount1KFaTILbRoPJXttbb0Y0SK9YeuaYe2LJP3BwzwzCtCrlbZkmB+mI05lxDWa
CwvSZE/D6cKrLowP5oYPtUcOXrQlDEIcRLvH5bzmkPaa6CILa3W5H1E4PdGoU4on
W17LKFMtCp4okY/h52lPCuLhnPZSYkBEAvC9XqYDCr9Cg/dMjxg3dPpa7ktVR1a9
3S9ZaOkuLeS64UvrQwA/wzEqGYxcMe9qMKeXrHSwE6FaVwgYVaafI1KN1LRWf21E
HPsDKQ+kaDeLodvmHETkoRUWSF+mZ+ABZnZjp0+jqzeCQBBSphVtEntlU7M5wVFD
BmPOkLmA0P1PoUs5oroAWSkzD42yva2hFt8hIhFqVHJMRSgEEACCvssNb3Axe9aQ
8aBNXEdGUXgZTiYCJzs2grDD975kfabw9eVVNFoEl0/jlCPgp7Odzh2rnhMoQspH
Jw556uDULDnSypi3GoxKsj5ZN2wh1GyZGXu6x1a9gs7+2gPMgExkYhXqtnboGigR
C4QqModgr1p/EY3s5rrqST8F1IZfOby+2/rkh4vGvHpipFBV+DuHAR9DSrcEI6iy
3Luqwr/8PmSUQ8KwdK7nZJNZaNRTZ86zup72WaNJnAeoeI3OOFk2A0bg/ZIM5RWw
LLgkJ9oHLlR46NaOr/+jBndmwUfYevAdkNJ+jK7oE/YXQJIjTt7pWaNTyiZPsVhF
7Y2enaSy9qnAZz5A/cfADNZawEf+U4VIuRWUWQizUeYNr7dCSN5zWeAudWqy378r
/CxGhu1i8W6C7nVDGviN/a9v9FkZiHhFNus1Av7ttnuT3KOFBiZF2jSBzWHnmpvR
h7huzvjSsCJSkdUArIC1iChlb/yU3e0Gd4W4KUNfyER06f4ludQzCbRPZ3tbxgyN
+3MAY/c1OrP41TYSqurPTrbvM8Epd266MiKv9Gq8dvIjeuQgSM6cctdqqVoBcILo
PaNOs6DY5MJqawzVhQg/rrDzHwdF1Nb+jLbuuB5nCeJ0Y8HSpQD3DhosorHTPUdc
KQbMmksuMWXFQym5BDjO+mX9h5Vj8Dlxo3z/wMwE8nUQUQqX2Dl+bdz9RwvKpfQV
YCjfxxjjgH+TZUxmtCqqrUQs4+RfY5WspPobPY50rkNSothcGbGcE7bes0dZe7tN
Cx94TXMe0ccSSCYV2SdX5+NLraDxxYB6+3YGH4wBbZHp6f65Af5RbZKnZLf52kPG
yBPVNbwp9tU8tfU2ZADf7Ej3aeYKiX42+J5E7ijcgnJ7OEXj5NiWb3eQgWPWLXOB
gIZUw7zr1U51GTsEo44hF593es5qvsoUPQiTQgNewHOfMT266fL2NZumHZHUxuvr
OEGF7qbaNTyOdvZFyHC9iLyyQgC1RCsRLRIOOYvIc3apCBtQ9YOQIBxYON1ecVPI
BaumOdZ8Ume8x/lCHBqFQ6dXfCqaT4ZpaApm/5XJrmzymwVx7q+0+te2hfh44Yzg
P5xnNvyBH7hvsxuACuFjckCrbzVGMdYf4Kp9gPkrELVuHMl7zvEDER3ZpsGj4UKQ
MiE27VPiemCOo64nCsprnJ64HED8elLgZUHDbWav4ZdLrnyI+oNw77RQxayqo1oK
vfDFA9iy2rUCNCZ3JGpmKRt6UlnAO7KaBfW88teOTh42E0lm4eTy2/wIyjng3V0O
OknMHUr61uzhfLOwg6xi40is80/ydwFhpS2uCmVwOz9LQMGKCnk/m3LgK1NhzpXr
xdgIsxRQbsZL9tLiwTTYBcujYmW6jFIm/Qm1nYS+lPknY1ClHz48beudyY+1SXcH
HNbl3x4hWIqm814JhNwu42V+pK4jwzP7oZnogLCcK7fdSpTRn2oHXzAP70zCxqUe
U73lfcVG/xWCYDG7wFI/BKdJgaZ+nYnC4j9ykrBzTf03q4w/Y6vl6jcJCfHT50WF
GefV/+cz5Cw2f0yQZ7EocF36YL6gRpqHEbEyldP4t/sIztJwHc15O8fItoASJPgu
ZzmGZra0VUTCiUitHZSf9FDA2OccRGK7mD1XdqGF2VJ01AHM2bwAgMGZsVK5GLWy
AKaCeycIstmhhRGW2r/1waRlgLdF2mobt5Wr8ZFoC53qx1Gf/8f9Hqgs+5QLVePp
vSVs/j9TEof2cWHEArpVkpK60YSolmcYNMj9HyPnzTunrXVA5cxxbYwRIeCOm/od
4Kif2iITbY+gI+BzSBp5motodNXD17FWAe8xcJWwkMFbWEdOcqOlK7FvqzsIA97C
QJ9/iF4n/tZH1IbTpfHd4PlRYiCpw4D60d7GvUa5A3p7vFmnPokWaeQxUC60qFrq
ZSmYH7VmdmjbW+B5mFEFJgoLue15zSugGDlHn5NihsCEU68i/5Pj/xaStlltAOCf
MnIWYxCvb2KGePSMlKm2AGgV0xHVGpdcowl6xoAoQzCEjCcO4mbrgS85oTGscgj1
mSI158p5nvW642sAwWWndWEeQla9al4GwmXOozWq7KGgEepYVTn97AuPpUmstAHd
ZjiqYVFdj6CAKKBPGpJdULr3qcBWj/VnQ8HATbfUEedQCmCLL3AYYm5cf00abJhI
jJ6bo1fgNInanAXJa2TPyCqSVGsdlXSq1VEAvKfT0CTtf0zm3Rnr/TYxHx6VD7lq
M7JXD5rImumhY3accYvhLwgQdoyKTH205f1vb3suyZ6Ffue6dRFrqa/uCSBB+W1Q
g2h2DAzg98dM9Qo0qmVbx5/TMJpmOdce4gHp8Kq4c1yDJEONumXKsNpnP0iTJp6D
Jv7Dnin+ctHOV++gPIPfx+ozEPjKZVoRd1XH1k3hCx8naXn7utQ+1g6K94fQxxfJ
aNVc3MW4jx/2y2mg53KgwLZnAonMKpjjGQLzvR5v8UDEr5xbjx8hy6KDjErQMc61
mLEo1Ja3nNP8BdUIltQXrboVFR/53wzk47QmB+DREFkIFTc56EyZ1QNn7kG0QvVK
5ZZnHf0HdQYrwHFYpTtqB1tkdnM5mZNAsNAk2QwsscW8DyFI2/kNf7CzDJujUZIS
0iV+TghOAXFBU7/ahQmNvwRkRqNhUD7wWM/6NSdXAqUEf89lYcLiayOL2u2VYiGl
4Rey5lHqOrBpRUlIpVZ2WacKPlRzT3CJDor1Y/KO6phveY2OeS1a2pw8OXF1zvpv
BozkOZx9rrFRR+yD/npWw8MmPsNWFWVmqnmO/lACOpFYkw25vj/dX59qJYABwFPJ
E4aIxdxXAqOGi8dpb56wdQGTVbvjkSFsL9Q6DWSC3ehThrm3THzMY2hv+/8aYtvH
2jqu0zjK+LDFyzcqpGqv/PQ6oBhu/wVdytdc5dqN5T84N0LghJj1bE2DJaaLbJqA
/MBsVskTZLjLnYxwSQusO5y4wewrtntHri0YsL0e3/wpVMNbZol52arFTLBiDF0K
`protect END_PROTECTED
