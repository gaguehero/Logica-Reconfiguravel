`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DID3drkhaWbtt3nPHRSEjxGnpLP9+X2FLowMwe2NvoB17zrj8wsJokg5LyKSQTJ
Q4ewKR5bJdZTV8LqyTKnfsU8GDDAmXA2bGxGt6GTYK1LloFo6dz5TX6Lnos7L3oS
SfT0UutY2ClPVsnLKddVejdcNFMcsDYQu1i9xqP6Y9veDxzVIog4N6F4m1A/dSwY
a9r4kLd2ER+kuHp2tasXcdptRf+vtQSmkrmwNpJ5XkWfb0gubHAb2MxtWtaDKsoP
DRjbzAUfZf4Gy+MqxoRqq/a1HGzk4MK4d4ZKAuDWir0YVXXqrKb7YHZSCM85yM3c
+LKA43UJg/NUyOIxn29DiJvWF177+ri/ioPV9XpuU+gNCrk4uzNK71PemNjAN06K
f2Jrnwv1A81b+/2Bo0nCpM82pVuexUApooMSvhZXSAMS/obaVO3LAd0f2KVdC8We
+cARThapQgrQGC9gaoWhAS+J/+90xXK7fBgRA+yGk8e35KP3T7K/2samrk7tG+Rq
ocXOgh3RyvwacV/1E/v4+ezTmPRVRpCgV3Qp2P4N3tiL8is0eKWZJnFJHfNJAEPC
WBps+FtQ81ma2uHV9gyDSZyeID2VcxaFq66zC2RxvmA185gqKD4bF0tFs/cboZHj
FLcKF2I0cKtQq6lmw0PzIcDdVkpmj1u0g12NI76eV6CZFz1X4ucE4fLo5i2PElaE
VbBxR7XFKXHY4+lznHwhWMcbSn5bLmd8K9YrDsD25oc=
`protect END_PROTECTED
