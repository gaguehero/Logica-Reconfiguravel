`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RFComBgiO5kAa70ZfiK3HUEkIQ2wNNwnGGy7P8YhEwQdm0fOUIb2HRwDtB+rxjTb
+OtkDgWiexEc6lDlTWBQqf8at+W2IVUoYPHPI+U3vSd/IR7u5CY0SFrukc2pkk4a
U04jlHcqWm66nsoSaB7Qxgce2Am1Qi02vbXwYWJxbNO85nfFIb9YN77b/92Pe1wN
XZNKc0X7GbN3wcMsEoVNhJt0YWbi6EQ8OZXkTuQ5oBU/EyQgneMIqRKhO2LZ2+tp
nFKxIQCxckZpWGdcH4XzB5AKKnAgSrj6zUFuhQ7QVYPW5H1w1NbyvGV4MJ9zM8XB
bgauPzgZREnEqMk3olIV1I5RknyVyINbENPhESo5vB2rHXtW4SqONqcrNM3SiGKi
maIfxwqgs4q8c8oL6npWpJ8kFSCLqVe1vx3iBg0cHMvX6grmFcxt/SRejlKRd+H9
rrM6C//BDwzQiToaF7PfMkHLEzPvCTRdwDBVj9hfJ1dlqdabk/hMbjdRimu66+hV
bixn4Er0Xe6NaRTpqu2w4SfhGSqKdGoSoUCH+H2kxoU3yiS1CBl95ZG/DEbhgHkY
PaGoaU/melN92QJYW87vx1s/Sa+FCbeL/jrqxMYqOkTTxpIO0ZF84CXi8lyLDTPW
OC7NJk3MgV8jBo1e7ses+Hv6qArQXW8j83CncACWcdqPo/dMS3Zf8G8fBdY3Tmj4
aOSa4MdIs+xAU9lvCvTNv42/eSfZK1QMkbAcl4DNSG5cMP6KFm2FXhNQGadTuh/I
MT7yi3Hqg2xvf9XMFBocQUPAT6hVGcTwPJXx03gkWpjkxiEZ1X+F+M3mFg0qrEIK
o1S0M+yxyYn2rtUDhWV06H+EJwrMkD/wEg9Foi2Apd8L+QlFJ/B62RYgjO+H8pfR
t5kC/ReNPVNRcIis9qq+gUC95RGpdXtoGL1wGJBBTAKbp2UGotcqhXxSoi6p59Ky
urq7XeG2jliYosfJCr0vqephPpbF4xRaIjnbBSdYtMaMwxid3Tc53ZNtx9AfQqDT
TRgtd2s50EuBL+yhKn0a/V0Z6jNDpMCEU6POMS78VPWLoMpOhVlzW5idGTDjBccO
KJ3qNcu4Wj992mqTDrC2lr25uktMD87dpaCGCymVy0SJlPXGHSUFqiKpJxushmTV
zzWAYSlzoP4BqLGAph/z7mQ8NxRO2qW5bnqQnD5kDY+AYhxefuL87Lt/W4KaV+4L
nwVlKuEuczaQny5F+B9eHwvGZvyLz57eVK2k8XjfaaiDgqnbnJcarqjKDH4KTQNL
GfZedRcwfs7r9ZKxEKutTqjMHhCPOI1sVsxbtMjmbVSMUnwpxeHyPe/AdAhfOSDa
AttAoD8qcf2V2630E8vy4/5124KfLksIv6AZXLtj19tfV4OPsg0sGts3JuLH+mOD
xh5U5B4S5ZXdC8rCaa+WlQi9qbp057X7WDPk4rHkInY5k8THHbxwkCTDliTUfoVf
tj/FY5t1g1Qr5kNVoPtEZUCD1dBZR4aBuUQkjxgS/tc6ws8h/2WcRA3FaORMsw+2
pqxjKLQAArSRwfNebou5u6fn2z28dkEsmJfc1Adpznn772XXBDRLQF/Mn41p733i
Saj/WffdKt+at0V8QWKoxRysoed4RFF6DwCAhwsi4Ugf+dSYdNYF5QbinnhXixGx
CWmgh2+NC5sItOYEi7+U9OW00+zu62lw2pZO7nHkbSAqdwifRGgac1GptFH7Ydsp
96wAXHa6pjx7yeAIHf3Eic65yrLe02hBP2jib5zTVxwc+EWqc8XQhBoIVKf3iY4c
Xj4AD0oj7Hh00Xd8hUsbUuIzKRCy599Ic3Y6rXaqHgpKIGqT5K6/TylqW4AINZ5C
HFV46KJKxYWV5DdPNuMDy0y41Rinn9YB+xcl2JSINIA3MIpoUDR40crLTKsE9GFB
Y7CusoKCDhQe2DouhYyzMZjdXFS1xu2H2Xq8jyW6iyHdD9ZnDDdWS6Cq1rRmNCvX
9NhIB2f9V/S6FwJOBCBDNH+mmFCefx08Q7cwmXcH1L5yWdwX4pePgiIFlLh2w9Jy
l9jQoz+2lk22xDN8Jpo1HRNLsb3OBnpSACH7EWoqtUsQdIz8o+yVanu+1dRKQBy+
CE74NA7m4EZshzNgc8/c0F4b5i8dVKA0AJ2fQ0YgNbfEw8DZYurQ1GtJ2DlVD7SB
pdzZ9PWwpZv2WbHvxlQtzH6qKKigWWMheuzE12t+U/eNeyJNOGv5dMo7xFBjF7lL
L97AnrwlTZusq5i+1FYujDXh1kfJlpc4DtDkZDU+TBoL7sePkiAfYlbt+FQfw1Dz
xi9D5dgy5i2aFIbUnEVb8nCo59EmbWGHnkHTqKaVWQc77iYPeQFE8SFEK7LaOh/r
Z2y2tKGuFGuG3f6YUnfbqLPFbRAKSFRmNf5pU6s1loc7UbohBy02mgKGiDKJJAZw
+oqO7sHOcZVySQu3d3cgXQbC10y4QkFn8hzz9X2ajinok/tNd96GJaIiU8yqsXXo
oOnZPNq006oaeiG0HlNNr3cBT9Hu/NA5Huwiv1mGnzZfWac+/H0LBOFqef6BVGuO
5IpGEn4pU2buWdeexhX3eqZ1/HDaND5aGnfqz+MAc15cOFCB8CUshM0SQ3Q2wB0l
eYR+X7vVmDLruma5+KNaTWUUAQHy9C6FKZwbQmuUzZiNHrdKd/Idt30mj3h/WsER
exYxTcWnz+W2LX9n2vMaRusO5DDFwclPWh1YiucNroyRo/hDYBOsW4k+Our24hZa
75wrkw7x1hSagQsIjEcoJijQpkV5YTBJQlbcm8Vqflv6Pw0BlviAXK6W7u+dbKu9
SASN4b7mtIAcisG5lbhYK9aFwDdQR0E5DiIQOg5HUodXdk/u2LSfrF/xreGlkSZh
BNL3PCBaMTc4gIEawP2Ud/UsNfL93xgDDq3EskHp4qMpQxefe7Wd2Ejtn4eY558/
DpNR2VmQ+RDwUt4fNmK5zPt5oFZK/GZCFJyBb3afiqnWthtmNy/O4H7I5H/ypPSJ
Fo7N1V9aMy7Hq1RAtVo20Xcv29bkT7OCZVCfw+ZIJpIYOpK1Lyr4mRvzDcZTpLuj
uFRTwqP/DWeF6YXQjLDplpXHIF/X75BwhV73MVLPfr66m5I7ApKQzng34QS0mCMC
I317M5zJnsAWJrdZmbMPs5Yvy997/Qq6WelKWXM+vbC1OWtcH8/jguGUYSVfP5sp
NdUXBa3g4G6MqAtRb0yJA54H20PK/RQadDKDGuB5PlDX7GJAxGIXLENyIfuZU5Qw
qPdPZm4J3TBhJ5x78gPTTPGNSSZMVpEzpzpvMF6rpA8BXgDUbBZrmY0cfQwtBulr
uU1eCdrq0ByaTCXrLKxen0Ai0FSAAfugod3PkXv1tUqgKSyS1ZHWoTdoc66X/H7e
5gT9TILPOKsLBwXyD2voPprL5oO/97r+sQ5BV13wknQqOiX3APEr9IbLmW0UtD8+
NVv+3IrCGemgy7gJj1NnGBauEOB82etZIrWgGXkv3+GebDrCtZDMNYNhrB28ZHmp
bLSuIkqqK3V4kCo46Hn0Jj9c9KfdONiIwP77KOU3XuIWEQo1jiEi/X5v7XBoxlJv
1STWtNQJHKm+0JI/t49K8efsGs5W2gRtEVXnrV2UHouIWrRNTOQ5syFtCPTwIfkW
9kScWCbr59K4FJ9xcJDkN+dIHdWXs6CLENcEyTK9UZqf2KGsiDIMoGOe49M1JbN2
7jjzffziOm8CtgNqPMSzmBF5/n6Zry9hTjt7OhYDYIeEbUPTdWjjsCY/c9Jqbsuv
LfQ8QMWgKdInO7toL5iB+4zjHzG8SktEF7N23OUfNScSTmmxVh9dAVSStb6zfrnm
+1Rj9ahNcoRPTPYqAMjKCQqMtv0VIro9laLfC32TwBd68peKBRH8BH+m5Bz8upFY
FDKLYOCBKclwAzN5mJQTH6VRhPNqnQvOg6Lv8s9Qc5Mf2lrLbVTgTHoRQNtxSJTB
Tft0oTxpecw2xr8uY+wJSCP4yoX7tULXmGED+thiJUOIQk3iYA+TiZheBNoQylEL
r0YeVCgga1pRxzRo6w1/4+kW4bSk4lcKhz8cW+Lcjy1IW8e14MhPx4nDmEQ+B8Yt
StTT4BdM4Zf/gmwgS3SDdQlj0hQ5cE3CrK9XlKpxFfuLBFG6tiyuZ0LspiYUSN1Y
IpnAF9NQQOL403PFC1xLFdqpMNchOeAFz7fCrdxOsI7JhTy8KeIDbWzdcrDHgxKN
Uj8vRPKSMqufinSCjb94P58qIt/5zC2ugO/fUPRYRCzdYYUkp82RfQTWVNS8KPcf
x4YLM8HAy4QXLmtSi/ZRLcEqTPEr0h/U8rI5AZOIdQwpiodFLMCFXDqbuSvUL1rb
4OWrRUDDhJjDals8YsEhCtHRl++H8DQJ9jLkOXWSBYQNIwOSSHEsw6sEUDMXYNc6
W9JfAUPb++lYsf3HWMUifhV2ZepKiuuVDMI1W02pppZPkjYrsnW9ZHEWhlVDtkHn
5j6YRrXW8ZTdovYd5E60ZQOHJa44q3qQhbQ4DzWMKnZ7pWVl3vPzoyt2gmeZ535t
/rOzCkL4Ro/RTk4boSmNn4LTmbDEMyaCoxCbHGGL53kIT4tCAno1s2AiLigB2tD4
Hr12N1NmEZMJ2Owlb1TRG9cfi/pKFGG6qxGiQud9kvog7vjvSG0/C3DWJv2lWajy
/xRjZ0dShobGa7DhL4WLtFkySco+CAF/hzAp7kuE1HLZitLSGU275YZ4haPSv9hL
ULOzXJmTnvbWkc+RzwvgCe3rWcBdEVdFXUv7Y39MhVK6inmXJRgKhazQQxgy+nt5
8mwoHH2XKBNou7qUc6gwojjvUS01RfDwYO0EzQRTv/lb+RLxgx/5BT5vTwgHx2AB
4om9ZMOsY52d/CPfGWc70MRLf7Bd9j10SRGQ2Ijl1yeiy9U19bw5UU2lfjo+zIkH
ATWcrEedEMGtEHbMdz9ewKXBQTYuN8PcdCkp4ksF0hIeVYqC2NupPrVK5C8oZ1/x
U02w9gHESlLlPLna/6900VwQD3jxMmyCQLyFPzKJWvs+IggBKEPKkykb1VpM56HG
KyieDk+2xwo4ChDIs0UFO0UkML8CuYMCN2azisRIMUOom5RiFFp7gtaxylc/AAof
xge8Ns46qfNsJpNivKCZpOEpZO0hdxWIFiaZ3jjZGUDQWO6WVneiNh2fJWBDKcZJ
597t8rtGTCoN8PPLHxdjMj5jv0rkP6BvNnxccWl31U2SA9Z8JL1/T+ZmrwlF/mcD
txT1POOYMCirX+c5ZyJw8mMn9jzPGiRD1zmfnoAYgAgvsFYakFaAGL3oTNs/4hHp
mGK49JhFpqVTrLNdUOTRWnNj71Up4jYzHmjohz8jif38StDZl5tkspcA1GDDa4XE
8e5jRejUR+Sjlb6NY93JleTXyYRwmyhcvqqU+no/Vg4nKXwn3nfI0sWo4mcGLF6B
m6NXb+glPi3UCngU+ypk6yBo/p1D0l9DcQ7sCm2qWyfGpL5yaJOtDux25bl8MhFn
Q5xsQMpdmKj4yqSz3srVycep/zosWEV1eMwXknzQ/FEdato4ldKkSOcD5FrnXtd+
+cFdhdF8PQcQ532/YXHew8qvysEvbtNTWCSp2LZ2TcD/FYHwMmaoc+Kmmmub+1PK
I2DCVBvfnKJJwtYkek4I2ODt+d1Dy0xZPDW7+Vnh0rY4fIeR5LS2B0s/q3QSz5Br
8KXEh3KhSjTb+Rx8Yr3WZHVvCiHqPsuyMeTC+dj5ApM28GG4cfsjq7ZgN+T5nPzX
aE917kVYXoA1tz1eMJCvaSZ9qgseA4FpccN5wAEBtJatWsi33oDXSz8oTCLRBwEH
wo4ypDaCClioauJqw0YnOEYWRZGP1SJ27FRtqvsFvwESKchUWEi/ip8+Wk3R2Io9
Ja70+PCEyuEeL3DmhWfc9Y/mSdRdwFObncBcwTc96rGOUpUhe0du56Gwtj+nbZzi
vBLV/bV9ia0QzarXO/AfKVn+CRdNR2Y6evsvjpxsoKwSNsjranAdtZ4IaL2rUpo/
QQ2ZTSmFtQRJzMgKEeRLW+4XXOIFHVRYjDP1UOxHwjwMXnUDFbbePIzZ6YUJHXZe
mF9F8ay8wmpDctFboA8LSH2DbSY0mJtg+Qvg0RtzhdwtLd16yR+IH7eYNbebZaui
1PN2BVR3EToCSpjY8KwIrhGwcFkwLrIUWhlEMrBAGsyvp3UyJKQ+L1nhIvq9f/Ba
07G6UXfuWPdbUbMWARW62t44JwLJVKPZXDGM9gKBLQfBx+B+pVBFb8vpUZoyXLdc
YJvKrLC8Yh/c1Qsjk4/GiCyQzazhhen5tFZMHS+wK2z5rNn0+W56/4DD1295wW7p
KHMFNPRZFGA3+3Rayr/U1/BwtXH1emsbjNoD9BcrjcQGA7UdS8tNVElH0DqPEiwE
+a/oyhCXhd29YdNoLk2GO87cQreMy/tvDtNLfvYHi3URz19L17nJ4DJTHqEMUSxj
UlLxjLNaoBNNNtRUPakWELZyaZ2EHUDpqHOTFJyb6680GPgGB92yOzQPG/UsMsDs
dPXnUuk/ZiPdgdrAnWbOcqx/13ScpmbXmMga+lhf690MrwZBqM1i8UBrZCIqdtmR
H8kVg5Rw2tOqc7rJ+3SRoMdBUfefCvaqzTCg1C3IwkcezOq29M9brLWNCMIjAOBq
/9JJinZydR1mO8CWJ62PF4K9IKUsKQa7hFoBo4WnJCy32GfYJy4AWqtFw/hy/+Ph
TlIzTFyk2441uq15zPailKUYMHMG1rYTJSc42DUgIUKT/ZCHGUmakrKix4xf8iIz
BshpEfTwkNCa3LnbuEYbsfLyfcl/lILrVJcSdEB8zwtISjm+bGTVJ3iZEaS/m/XY
iV6exPRMqMlQ/JuAE1DH1MgkmKo11eeMPuA4Ln+rV4EJJJCk/uVh0GWZ8pLpdUSW
Zht0FgquWzLjS2p8VmXQotzGypsrcQsAO+FEQrjJRNQNlBdZ9kCnJNBfk5YAZ7A1
VnxuzWYJyu3lFbKCN56bwALrlCYzp1qlnkok+xpgUf3JirMPqkp3hR7mSl97iugt
jJ+figxPBKRY43xYMOTCyVSFtFqhgk3EBZ9K3omMIXSGKDZkY6af0OgVKb+nFZlQ
IVqg4l0cAIZrKs0PUSDYTph5ZKYOpp4a1WjZOu8cwgoUGEkcJjvqwAEp/S6Nasuy
iE44vpDTXyef3F8CueSbjf9QQ2xyfQ5I29m72+z676bro7hB7SfnRgs9l33eQS0Z
bAiNzPkrHEviWJwILD10S3XyZW+aQEmKVe+7wHVBD/jYLJtUERCvwGvLYZLz9D6C
0h8p9rs+lUNpmQ1sL4u/n0So0B9ISEj2aJuFPTO4IUDY8WNklL7EvuwSyI9xByMn
7F/D7bbjA6fJ/h9z7ynCFc/vfH9bO+HACy8BkxZWBOBlAMYvlvsbnmC53zKC0Ak1
5Osn06x9AUvc8rgmOndIt/be3QZH0g8zCz657/pasXqaPyP/0tWDh5uRoGD+PDDs
9XCW63j1XTkBXJe9usCJIKxwcrbiDziOfMTEYAC9UIw4iuN9NyOj25Nzqjw6MYPc
Sjw/Dotd+Yn7gUWYNn4tZIh7ZjVcHP3sq9Y4KXGZaZdRxV9mvFJI99eWj7cHCSUW
yF5rSYvaBqEhNMbmeK6mAVW1qqG4eeb4GT/rI+W5Nbj32PsNCjDKtI2Jm2cfGMIM
`protect END_PROTECTED
