`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgWdKWi9Qz5BDyQ79A602NvuWEoLIkNz0ONE5zYNbaptojVuk6fXc8POSqdb/KuN
nvs+X9HpTLQddxJ7sejDoh1vMZ0XUD0Y/mf/95IDlZSxwkIha2fzFt6Y9kjBBcRe
2KnH/mXtT6Nj3n8IxF8mL3HDF5CwyIOmMV+WGZb5Fir2hW9TUd0SvqwyQ71rpPke
hFbfkjw1DCAwwSKioRuTOHS52Q1zQx+2bWn5wT/Da+O4b/GN3ZSK5i5voIR3LjPY
vydfTa8sx8QEe+8lot9u8b+ioMwUjRIp2x2TkYqpQOIHlPBNXexUyhPY5rkPdE2W
n5/fxK7EiJEDzI8SzrGiveM4zRm5lRrWJPtHEBxXsb4FhfprGAs54D5pIQJTK/lx
pM1cxFc4yj7Pfz1RdLRElGZTljdhcxDZQgw7E7x7b49yjNnPJ/ErQf5bv7O1tk/S
wf+7FNa8M6okIOUKVzihLUGWOpxAx5lUIguD4EAynf2nGoYr8pTIMpN690LhalMU
MuVF2DZ0cRBYlRpntYEt1NA1RYTzxiLMGhCkFfNkxh8wcMa9PkT0w/36D1hVygQD
w73w5yGrPFNXfol0bSvDi43z9yN+pbNYair/E6xGn15v6zzwSwFH+nkLC+MNx50h
ugfPyFlNbrnofUqjp/BN4yghiIei4Bcv1ejng9eY9bn98J1ZSbeR7FiXgjqwkfL6
PKSY3nlzOIEPe3Kw1ps+viEgL5Uo9dwsrvq0UX4xoEmCGhyTcBgyStF/2BlkFgae
5quKl/2shk2h921HP8FQTXOCTL9MMnHFgMpbu6V9BuTr+8+q4ooMOfY0dggT2I/S
SFQD8qOGZBw7c9hAmu4hkhz+ZnnLCC351QUaBMYMzP1aRsXDsYm+dRPv26w3gBGU
GOs8NrMXvHZpAcU4L8VWbXCUkhJ0kkEbVOEAZQLMzQ7RwcOKHlRYGsHKMy7BpkGS
fW2qjKEdZoTmLibS4x+y9KamdcHHfELcsbhaWQsuoAcQINCdcJ7IozQ1fpfUJELu
5Li3LlWWDy/E87WcdcWslw9y60Ql4m2qG3B7AEg9Vd558EttF6h+H4uWxnWWyVDd
P6s0dLZtbKCNjqiNZfA36CGCH8Cwsu2OLJA/zb2pSsA3oqb2pcCQkigjY/dtr4FM
BrV6lOW9v8G1uU+kE1iZB+zQfWPE2u4nlpzmhDiBE3ny6pQovCH8+szF1FYbBtTh
XjUnbh65bKADRFkwuideSpwGqwwpwR8mY4PXB/T6Syk=
`protect END_PROTECTED
