`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlPhBCorqPuiooI0HcN91Axw3lDe4TCRKv6I5SbDnf/CTX+t7a64fyvuf4MoNXOw
OjNdNme3HxhAcCJRDF/qFiXU/+Gpgmdw9g0ZdEY7MOtIp7F4tEh2vCfRj/OC2bEW
ey+gesWkdZ234k29y7D0vUuDHOXebdRMvw2/9F6W9s9/AF9E3TtGaxqkpA2fniCr
MTiXO6gxUPtgUYdTqYSkRdUicEAZ4B8Oe9FxZuL/heel70qWCfxaXJA/01QXLsW1
ze67hsepK6N1eGZ+lpblCGOz76c5ivSVZ2WK4ugejkRAPcpCNQpdm4MXJvmNE8ai
a7aTxs0l7DnM9h8Ry5piotYbocifUjeJSLIAGybIlatCunA4V1k27oxL8y9e4bbM
eRBCK8kK3BG2l6hG+UIa2C4y1GD0MsZFcc3gmpmQy5o+PHTynNRw2Devhj30reRn
Q/7PAMM2RZySMFZeGfIJ7Uv3hIbaMuXbMzqDEMQKuKqcYt06QOooI9UPKL4WSvdW
J5kaU8WrV068WUJ/7CCzXlc8EhoIo/e4L0a9uVTz69mykVEx1fE6CCEljp/LWEDR
DPbCnXFQCQpOtir6dyRX9I2SVK5bA4vlFbkr2OOZqCvffCn4tDhFF9Lwe6ikMtc2
eSvQB+axr6SZ78WwUX3STVgE2CcQ2fpfalRVLdl8TEhmo6MAhqjkOG+9iUpCQNSw
`protect END_PROTECTED
