`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YG8EN94hSxtlHjWj27qyo9xtHzdw6lWBWuOtrzueDj7ILW+XiQo/ld/LWCxnSAzy
MHDMm5agBM47G5AfVsqd2iRGlerZFfzz30H6ndzJ1hG5LFk9XnwqUHRY4KAMdIlX
iZM4gijBBoCAIrxaQc1iq2nfpnBXSMpxWRQPtGZbyb0MGFM0JkVv9JTtBARS4D3h
gMgDrF+oBpCr/vq5gpEzd1zKEHVJtJSGpPDmmN04rZRwg95xq23TZooYmqJdc/l1
8vWkEpKDkge17jUVaE0kNgUB1TNN+Eb6LhdwJDCYogUT/MSbaLYFv6UktHPMD0MN
GDaPZSPtJBgJmaIP6e2jpO6Ggry587z2bQ7bTzG8Ntm5Xq/e+4E4Tm6Hg7PebaAR
twOkV6cTs5fnRmgMf2RWVZnBkVSi0ZqRT704ApKc7FDf0YQOt52sAztH0/mXlXoQ
jz1qIyQkTlgG3OHKZHASgN6sft0lwg8As8x/vuC+idO3qx/OihflfOAbsLaMDmzv
j1akhvDYTL/V+zflD4gzjzirEuRItW6flE247ZgQI21XZfJVfLnwMljOuxJ6p8PP
w5xY1mis8X5r2GYOGsl50N/x7bVFt6y50y4sl0N4+/VXDZbIZZHLUybq/36h+vpo
jANUA4ot1emEkBRZJcH5V10ur5gy330tV6+sF7TYRfv8HvSmO4qb9w9HPQLAaVb/
oo7IsoZ4NmPWWTZzeNof7POFmhxG9irF+7KYM90RyqqTHlUAjv3hlv+AQ/pFVCTm
OJ3uhgLpQVNuj2SqJUyP/QIJPwH7p/fGQZuvX0JdtCsnRfILPnehcs8wWIxksY61
AJJw2eMugiswHApR60ye7j4V1lCDWs1JytNx4As00L6HUYZ6NITuZvNadoqRD6OM
UjwvSjrel28msVG5tZ0+/T0RKVxxC2/bf35mSGlU64xJwnWOL4cYJWq1jK4c6bI4
kMYHVKshGesMrnZZ8Q0QjR1QueSky4TnXO17Tizgqdsgjzw3kY05wARd7MXy+sgv
wyn2s/kuNU16qX1FtM39tPJYhCR5GZRXh519xqiLRJZfZ1XYNV4IDOmqGn4RYtp0
lw4ZwZ/y0rpfj9HwOIfk0ygGFhCjPTdBjag6Lw+VCuTeullMNOkZc8hNRwVlSoHJ
Qafpp5qbaLOpKG2t46RhWWj5jLfylrbZikYJZIqbQsl14kX+C+tyt2kdBM40SVsa
uCFj7NTCTvUtBOYyOZ0P6Q/G3iZgHAvCy7AxHgeEKLk7Dx2Pt3uejwg23VHcRKJZ
p9Rh7dVpwTseu6zRAmjnvgHckFlWXPlACPCSjPb97Vh77BZYwWec0GWvZVZNlSXh
/LtsW9ZyBTa8hsLTgnbJTSou9wT37GD1Ks3rCmtS+kAqD0e/rsSweTLS4j4TBmlY
VaQ2KHwcVmp1GLObrgZTqRIvT6eYuirzBopx6G+4k3ojCBHDc8rjX1pQ4iHQwwcY
VQDuZliOBJ3WTbnDSrQWNA6GoJgg7WQWA/NLGFcFuhWBWPQUmIgi8BAV96/7BV3n
XSwJWZuIwfS0fD8vgRsacF7JXmjM1Tw9TGXu+I9mNKENOkhhw0oJToleHjvXomyK
ouvZPwFXFPcpXlXXVb5ga3uy905FqDsTq81kCW+4h07WWBDveLI4vmGyYHLDagfE
+BDnc8/jMxi5EjSoarZS49lWVSH2ap7jYqR9b7tYXhUlFq4oGWY1wdf+CI+tZLMc
KbTtIVMkt97TDuRJzy7cXete0WiHY+X6T0JAp2eNAmXyL/ljlqBzM0kK9/qd93+d
lqlEqy7voVI4xgoPqe3toLKhRTF79khkolxCV0CTfIxyfuqyQIks6LBQWiuGs6+7
R+j3QJUAYA6FD27B5fuAEEUn+yo2x3TaqS6u4EkPXKBw+bjSITEEiJwWU5qGn4BB
L0Y3Twy52XaCykTFGpTGsOD6ofyKz68aZF0cudHl8XkOw3tbA5F0zZpPILVSd5Q+
Gg+7xWeLs8C/VF5qy5SsZWFH6NFR+8726o0226rxrxofOpotlSLOYfY/1KIZHONQ
`protect END_PROTECTED
