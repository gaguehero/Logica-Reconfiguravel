`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tF4hOqRmHmlP8/P32fYTv1vdZc9LILi2EPg8tucjKYD/t8aVaWUdyDJ0qNVwQMzK
aKso2o/qxWg441ceqq3ZJ+1+YynnDAf2zjir9NPKN2q4FGjt2r6zr3NMObyE7/WU
oEKVJ+h/8Rl/fkqDLUDkoJKWZeHQMiKPSceE7KTiulZBCtABBXJVj0kN/t18z6yy
dOp532hRcp6VgygFAOPCQte/pEblGFtX4Zisa3sHpv1R2dU4xG2x7lEhtuRl6Z2v
Rk4UyBW0Z1CQbcF61L78++hZwph8IYsvCRNPQXsGzxp2+DqRmfzS1BC+jrOY20rg
LJ97wb7Admbcp+WDiC92XDrZw+lGBH+/7OpIoxn49fo42/43Kaltvqy6OHoEXzZJ
31sr/zXwRyHeSxyZEwc1rOyVtZoYW9PugBaENwJnC8AAwyqHVnbOrOixP2ex+nlX
o+K3bwVjaik+FSXdz/KPRmo4uULMLIwAcf2NG+He2gZ1rwfhkw+17ls4FsCF27YH
Fh9VoinSsgB9ZRRdzPeHQEN1KhW3P2cqOhPot0s2kxtRV4IOCWC8AS7QthhhjZIh
uJ836oE1wo6+/sSIswvvp23PYAvBIIkQULaDDbUXbrWVQf3nZLQclp7vRsImQwZQ
WmOWRredseb96pKTtjFwSQ==
`protect END_PROTECTED
