`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7QFFxzcMdiEQUIqVEtAF/6Rv74BE7mmROGZqCKFL6Hft/QtcVecTtoP0otiHERd
fDMs0l6OkuVbeFhp+RlemCgMJ4EgTR1mQNtqoGY/vyIPi2BnhpamcjK/H03t8PyM
2J2Y+aW3bYi3X6pWyb2kbJvyV77eNWM1gpurJQ2UYXrq8gS0R9leWWrBfap0cf4m
IgdQJKVA9VNAprXbruMtwCe3k1lr2yQgrWHqfi1djBicATSPYFNC1HOZEShKgoK4
P4ks87yjTg5dWaGwolErUljpehbzNpPmYsM9WdvUSMojw/UnhFkxJEmmLoEYweZO
8NdwrbD+8PJP5grzeaAn4alo5kTSxO+vzpz2bK5Ecda3LF2Mf0tq1qgAgPa59gcl
v6M4te2KHFx64SYJk7fAS4cSbT7tf1PbrRO0qJiPGCRtjAUjh2cFDoRV/6VW96mm
oJ9ddVCxeptbwde7NeXO9DClHYf0iU5jlruG3omqvcxY/7MqQ7NhmmLtUlTari3b
XOMiXK99mTXascMqpQ2mEzwMTaUrDIiQxY8ctUEjhHm1/G4CEjappQnuaxryZ3UY
KZWbGTKs/nMqUvcIfDfgRyybHM+avDpI7rTfFpJj7s3vfj9KcCK2GiJypETEYlqw
4OrQcrIowfEOxI1/ffhlpvSCIvvlVy59pVhYE6jqzVElC5tYArIsv0QPaU4U29lP
wlMMq1t+ottjfolH631yN8vj+/b98ewbMpdh5Fz+xR8kbuPMjDR+l7/7UPYWVvV1
yU6Ib4HMuLrpWo0ENQ31sE0QvWepEb4IkqvX3+Etyc3GmCI8+R9F6C0lLd0FjS/S
4bCv/5fzQFKFVkV4R49NrFcwgkjOyiDRT3A3bnx/753NDYZhXmhGBJ7XshpDIQe/
R7Z2gugZFR7HqLHPG0aRuXGN/68+KjZZ68wU5Pa4eOEFIqawLi7r0kjVj+Wj98eL
BqodkEF35QSkMKmIxmGmSoY3yT2xBNgPzqC5eJVtgM7puhOqfL1zMitahX8cB/sO
1xJ+L+dCcklajM+FRBAMcP0yaNPrc+lG6xatkuUZEo9umZxGYHaH/rDODu0JtLZb
cDO1FSndnIkT96a8ykxsQoyuDjnPzVgXjwnnX0PXtpOgE5wEV3IOWxhxp1eBPkIB
DnESpknv90lqPKFYI8lRpeFSWo3lF+0rW+Q6Ud35+IYI+kLmnW/bV3HlfBLdOIut
NVf+diJCl2VF+KIcViCGRgCzimgvavD/FiFnat/EZA5xYAUG4MDVibQnVgqYni6q
ZFfGHS+9PuC8skAvXuH8e9p27WK6up4l85DBlyPREjBzdXNjv31wp48OJbY4mKUY
3SdUFCRd4GLIUbDyi4s+Ktm1ilvxNtREWplCjh5Xf1ZWj79mmOQcbMPAz8JXf5Y9
9tCrdO+LVghwVb3CYmCt4+dtyFaiVQMWLes1MWMxwmBTrhbHbYExQc4uquGcUqLP
Zht/e/IGL2MJBkmWosMPjM7nihEIfif3WArYWUGZD4L+R65rm+j9uRJVGdeHk1jz
JFqZyyZtOb8+jByRt0VgMGRNp9dBcGi4VJOAlZ6zCj1PDgKyhK6ZcDo6XGyboiRV
am1sJCsqP1QCU9zSXGNudBXGMmmOTog9N/cmmD7A1jzxvdklCvpxy78F2tizjoS9
r6ZwgJOoeKOmBZyASVlrOvAWwh/gUcn93+rBP7jgbg5Dt+huiYvZAvHVGrYdu4RE
/I1nrQdMan08kHHmKFAO3QXfldIo5ZDE/Xnh0lFomiXoBB+y/kAY19sfiGKkAyYb
BL7ubFkmmb/d4qpbC8FhSl+UAh+COm2sElbQJVerZ1jEPVkC9mYOYyNtJhlVzPvU
IWNx3PQmnm8lZX4vPMjVDjeOu0d6hVnRLX42uEIrJAAcyBwu+99L9dWJ/08AIzfL
vagtFt/YWf4+w91jJS21kftc4EM9ol5EYeYNcnxRtDIBT+gqXalwkRtGOdIMNeck
2Wa+D2Q56YqBmoC3YnlVMnBzQCYfscLdNdH8Yss7xXS/Wrl7ijjh0W7wUNV5t4lb
`protect END_PROTECTED
