`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzQwEumUnuDMMOX0tUTrcUhz/9fPjke2fslDCpsLgaRaeuUTPFXGfVHis5gf2ENY
fJrqSOGn/YJ8ckbfkSYrD1TLTBcSiVu30Te261aDgsSDOoiUH4D0bv9IzbzYXaDX
tMjx5S+cyKMQd5bzBUEXSR1KRPKl+5ba+m2LyZRGIZVrRGQ09uY4vPNkqBLVMkFv
4joPVUCz91LiRdD3yGIqmg0Gg/GHnkDMJw6gYUDMza0UofDSD/mb/Y/xvqxRUtL7
n2azN3SN+51asOTaF9lQL4Aa/RdRbAKPS0tBV/lIU7T/m2EIS20Rc0Dwx8SWVkxb
j2futaJO6L7XEUzHlKhG0J3IkoyRnHvv4UJkxLHB6+b+q3RjaxeAiNYl6OQinSFN
xG1O8LwOjchcAEI3ARWY/g65wfjORenr025C87iIZSHulrSw4mdVZeR58nqOD/8E
Wm/kdJabzQwtxtUE27c0r1PqsdbA7NPoXQJk/Vh17vLK6I1wY44j9kNCcUyDRZfb
ZTakwWo6nwq7Ivl1DeIXyosNfAMz2vbTwehLW+/6a6Z0Ei8aVFWWNjC0utB1OvwI
yRbp5b2q7H/vkZUkJ9dD8KAPb/hUgpbBaRnz+5ykUUIG34s+pykUHOh/83vnmyR4
aTWH+iSzsVvRt7zmwB52EA==
`protect END_PROTECTED
