`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vf+X0UPMYXFxgW+bLUooGgbACkXK/WstANX/YWciypyNwNhrtJ092JtW0J13QzPz
dTwdu1Vabku9mRvPnW3fsW6XI5kbD8iZVWvHe1n0AWLqZh/Yk5GiujfRtd4hnu1W
bBy4ePygpR5vEryG0/eFsyR+8JdT0sr4fyRUmxkcREwctxx5v/MeUqBVyB1HUoV1
G3wpskRVzt/aADIeUOPl6YP95vrjMkEHvCR4HvUqDY1zn1uxeGb3Ik7Q2aMSzy2Y
XKojGvMkyHRz4+j/mbk2ep9fNS6etyF5pt0QfNU6iQ4OW4RPho39zBKo6+CWkCp4
bTvp+ruVBC5Mpc/4CvJYNEsJFGkRdEmOgegszkUwfjNa2lonz8jG98YWZZb4koGF
bSrOSSE/3WEuuChjgvA5L2bV+fVa7ysbppjet0AXSlI7v7qsOeplIovJy9+EOcO2
bd2JDRHct87aeh8gnE6xyY/4Cd45Rb8b6cv2QGFUV/SolYlmhfRB6GvSL8nwA/8Q
KKghUA/Q2ZOd1UTCE0Z41eu2Pgd+zOWxqYiGr4aboRWpg5Bu6KNRneU7WJMp3pOm
Sad7R5iwDZ0mXWbr46X2TRUsFDV/iJ8jOxZjHznx3Ea/fDsHdm+6IhkUPZsx2fME
jcLqs8Wqv5j7xV90pHLWAZCtx7hjheRTVJq9K1STcukXPCvIDLuSA8X3X4NDAxlY
8ut8PMJZoI7fkvYh/vN383FmKctZHGL4nWzJbdH97X8=
`protect END_PROTECTED
