`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WH9/jCbDV0LgV1cAl2p0qhmrPS1tMSwHpbZ5PUJxICOkx4JNcCd1mxFo2Xjquv8u
q8lXbXOtd9A6FRdS2W4xkhMmYkzAF9gU0n1j1kqfzkkxeLEtOKNp9V3RHTl4B5zS
6b84CsKlemK6uFahcHqkfhNlnJrJaob9QIALai8DUl+M7K9TvJHgzgsTIJ4DdI9C
Tuv55MkJa+xUKmLH3vyc/Cp7Fos4N1WGv7Nx8ICUyPrY0y6LExNBTTiIHoAUKB2L
nZYD8x5jB6J3zF1eeWuFtnwnX+C1ztgmbrr3EIM51fbmDVDuqcgBF9aluTWRq5Fb
ugqjcJOYZnTiGMJJJhq4+0Tu7WzEsT7v3F5xCEFKQMvTv5h+wQPa8cWP9papkn+S
LquliaP6CSxGnjDFFSR3AfYMfdPvQhBxBnKUNP9onktpd6yIU/ZzEzCh8Ji1qDhb
t0RVMo9WqdePbXcgzIBaqJYcZZkEYjQ3ilupid8UXF79efqW20UCh6g549dc8Lq7
jRYSX+uosjHdWvcUHf5UTMkqZ205MB+ANnSkgz6JPDyzVpNlkrR1Vq11AIZwEJdW
c5qveDKX+Eo1M6Chn9NKXZ8gbAYUb6bhAQTxsdSw2SWmEGd7n+pPP7ZEVOrSL4a5
GC+gAk0t5L7QBcBMgXjSs2qJ8uUQ7V5l0Zr26ldmEnuJHB0gpLSqDf4LgBj0JYqx
IJuBrLPNyx7qkhG0W7fRhvCM5wRt8KHQG1dxaYw0hWAv6UP5GXGMNOOYcUfsr4rq
ct+MhQiF2Duco11K8xwPfMuwoLGXCrI2LAsIJORGjw4aueMuiduZhVJ1hLEIro2r
zI16CpKMMwVcatKTXw3sI0jwKE5LYRhoW+mDFCTteo3DnmW+osI3CWzI8QUNtP3h
B1rnS3o0X1dvLLUbH84JlFzVEUcGskiEiBXrFhWpa3ldBp65ln7iMmKRhtRq2ssC
kw1xn9Ufv1UVN+asojeSHk/KGQIRMoXgmHhoY2pFzssUKbNz+q3JyMZbtphs1I9X
n/zi/QM/os7VzZ8ttAwPVDsNuTcrWMJR/dVYD/P3QwVz9IJ0XbvJyZ5HFpMwrXUk
hyPQywkdzXdRSpkkFVeV3IGkv8F4ehQTwd+1SaDOChnTII4PFoHFAHIjbpSgUloJ
gxVw/SeM8Dcet/aRFDMjSqYxOPUJ2cumyicXmB8OldngDsthVadPtCAwpagIokL1
cXGeJZf8d8KQfH82jQpeBNbLiFAsStLbnuYIhTWYCOiXC76ipevYwEldvkAyF12k
/i8Wr8fK1rjTjWMfpEutqVQmSk5ZmbZRZQ1S4syfFR3jaF+Dh49z1aKS34lotr6b
7+q4csV3tWaxRLbUj4SDf7dFIo3xcohjiJK2iu+opCjveVbgiO7xsrXbJQ2GeFeG
VaSEGvbPVQYLWM3Azm2kRe0gm6wajdJtxVP7LIGGVHnF3YMuNAUpj9EyNLVtYFsC
KbwytP9WoYtHSp8l/O7goNLz0FeRR4+g9Py6UX1Jn74OoI5acShRD+XFU1RnjKG5
vyPjPAt4LlTahtqeLWhP6LZslmZDZrk0NOYsnDcssQsSQ8sr2fwCK8TysFtFfL6M
/WmQ4ikI/8+bN0FpaalugFYAXWJ2M269hqqxkdbaVg/Is1PRVi0VwTtRPKALJcdz
1B6FH/e9Yp79mz1TuNR2OYehJ6TRPqhI5FNqhiAcX7fLsFQlUkzloDmOILjUBiWy
RgZ47pfp0OK4TLCb0wUOWKsX6kD6r7RPRPNJzZI78XHGNu2SqD1I1i9CR0Z+IdA+
R7WTqVJZz73CQ96ffOCrApdcCPBfDOtCAHmRTiuN6YPaqOhKvQdfERscvXxv8eX2
4IB1UrSSCGzQ6P7hIlkMf8S3wDA96djI3InSzprJ7zRFYu/rY1WnrGozEww2GZtc
VT6NYekZbdDJe0Q0DBJcQ75vBQwSA/XKvoBtamzdPH6BfgnQ+rBZofMkK9+5J3hr
ezF2JrEsU06p4bQ6QPu3CZI8PHgVkFeSKFyO4tFJAB+Gu8c30QMAVf2Hj81uIfJF
oOLOFKISBj+gWx8YNIyI42iFSK5yZNVKHWgdRK6r1COcyHgXO0sw6Bs4wxNOKdhh
/cW4qPsfHban8d5zqipFLMRc45VlN4z6EDdnCIvC4ERheZOl5/Igfpje1cHYOnB1
ubXVGsUF2+CLHplwKV3ow8+Kgdpe7oWc2yIJmqCxSXe7wp37qJq1AG7EW/se1cw8
dulPV2HaUtAeSpMRtnYxC2FPyG93P3QxWvLIs8kozvpqijEXQuBOmZ1mYIAvF3SL
PVE8HgVhguxGlJ0NzTVWBwTuHWX/lqKh7CfTMSTaLzA1t/2ZEOM/gGW+Jy1IvMq2
0e8GhFd8ule18BZE+lwQvLrsvUmG7vaQu7WQyj6NXHgaIFJz3QLfj7OnXjwyTwwN
5nilWAWkpya2Zz0hAAWT2mIwetyswIq5y6GVu76e2NXGWHFklwv//vZcIKbzsBXF
CJ889QfcramTL+NlJYIbwweTaK8mCWH3im7SqnBeeLyvs3pKkJs5bQNaUqzpSZN5
rEwQuvsVgY9JL/qLCiWKkzP72lnChchH4+2JFmi8EJtqFhDxDwvChp1u28qW4YsM
ELC3seK4IuP7Pl8FqLJWuYC8c+fVdDeuqaQjL9u8qwIb01TG/CP1D9/H5gEBR+Vm
QjqAvx7LcLWMxOoKwj7foihxjfMrB+nCgHB2HAehYWRsOydIc4IIREkQq4A0NSB8
8MCX98SuvdgipSIIE9uxL4tpOG5n5UxyRzwjn+IVMrJQJZnHCLAr8+KtFpDBleIY
4p2TlfFP+dzVHk55eKW5vgrh3STPivmBs43y/KhHQtPNhC6eVj4oogNL5au2nDlR
8xWFD9YJahLgvvdPeYPiR5HxLCPJM1u0ToTMFKI/SNal502HfKbOPiCyE7vkzEkV
9fL4zmoa55FibP3CHvLwZ4IOEYSuwYuuBe/b0uhB7eVWm0vwFmWmJTlB/QuwJY3R
BUmFc3c5OBu5HE+e9Ve4gjHKwRuNZ8NAl3VTJ35xmufsQw5S+9SFMY9oJp3QK+5p
AZozlT9rIAo6uJvoZDMEYklFb5gFW8Rh/joI5Un02fxsaZTDVaUaU60FWAGI77n3
Vzyb8PLOQRWWff/Zw+Pkj7nk+lCeZSGsafUCjIoMQeMTzH0lVIvvoqn1KkMr2rWi
dc6mRWjtJdUruvVWTrJgF56WcWoKSAJO5grhRw7NzxvDmqOtV8dip25DZg6hX9m2
m+E+eEviyeHz5lFdE+lN1mLTiOPmn5twu3PqodVG4Y7mfho4HBbHeqhZYTGauDce
kLuESRmhUAH8ccGjgVVJ9E1bZjg8GKeKmGBH4B0oyjo7sLoe+gvCUv9CFBh/uhgd
z1MSM6wipX80FGLggUM+0RDKnmuH1qX8b5kZA0b1RA/zqGiUjUDDO8Xm2rB3Qg4N
hQX6HzTkkFL+HnQ09PDD/kdosT8R3GWlPnxvWG75VzzvHKTjXoPAbQmj+MfjiALE
xbDloL+9ffe/qyye72DJdLQoYk81/QmztnW46BNA0750z49HLLrcsP9dOkjqXKj+
Mpl1GkBdmVsT2974DKU2amtwOpdgSQfVs8RlDjhdUxNnBNKt0RWizKHihbLir+7U
bgDuf25uXuoHOUz2CdvuKWFloM+4tTFVPESEua1ga13mgMlYLRsJh/WaYhO88Dfu
XBg95+JPjXGJw98pon3hBU3Zql0uiouLwdFomIDqVNC5JGleMqXK69SOXbtt81CS
DOwY6+EI+FUmXVqBMb8TKOgVcMuNh7g6ndq5T57I2oddZWX36dDkvdO9XgU080+r
6Y3HzfknXsMqNrw/UCpYiZMjNwRmUYLberpta6KAnhcM/lo2C36M0nCPvL7ROTKP
bJFAt5tXmUn+XSh5V/8l+7w+CbTcmkTU2yQ2icedXsqqNAeg/N8bgFrDjJCxrNkP
ASd1pGtt5BnPgVEMHlgbf9/D0SMsStnOcGJmeRDLdRJx4njTq+gKsl4AXk+eg0GO
VVf+6gQbQesbVMbFGl/iJB2rtoFxNTTquWx8LbS+s+beoUBLKOdyDMcHzG0b2ZlS
Mdok/9UhSPOK3XR9Kf6JihgyCvTkRBcEaV/J8yS17bWE5Ikd5LPKIHxaBdqKC3NH
pyk7t2Oc4o/VuQRN2XBjMRoR8+vcSMFyoHllLbJj1fn/Afox8XOb6mAO45g0KtJK
1HLiSKsK0aq9kSRWNzOo0lPxbaLh6Ib+cDWaq53aqHbsQYfIGdUwPZH1c0SNv96D
7lzi3oDoODHMCW0v1+7zGYJvdpf1fNlqUm2YReaAM/18oGijKXuYkMrJy/axS9j9
Trser9VVT8YibmMHPwvVaTmO9Ga3rC1nkPfcGrWq+87+m+m3aK3l/nRkf8QmhsVf
BmFjCyUKnb7/0w6QLb+E7AWFYgmNt/Y1hFftziElI9ZVmg7qhRVAZ+CUOHUfOkh0
n54driPX5teOFq/ixOeeV1OSrO1Qt4xpLkyDusd2a1E4BzdGLjQp0swLS7hwEAc/
ehsTmW4FCnD1DiW7GBY14rP6v0cMaVavuVONJPJx2e+ISuOfmApT6/mIaEaWtVOQ
UA34edMpw2YoKDHz6v2gTp3x7Sm1/AZX3S9tbNikCvo8gVec/Lqc7lPP8YlE4l9H
XJP8lchob3W6TOQ3g282IOaAlGL9nSC4tyMi4ttlqUiXoC/dj96sRfuKdSpwglr1
f3QdwvxGh7+yK2hbhLQ+Y+E4heXNTRHVLeE5FTEkbaoht4PDtTCv5pnQVfrzAMuD
2HwGfI3bor0miDkrEnOeiwjMaitIWfF8QfHeSsdI7WBLW7S7CaOSSNKgCF5aiaOO
qsVmWOVDuzv/zMUvArNGngt8j+7p13DuOxF2ADs4aNgMpnwBvwapzdrO3snb2Su6
lg/XJsb2elOwPSsmpPaX0khfb9TWsLvCCsdyqR3MILC6MuLxgSLaBeHZQw0YETVf
Np38F+6o3/8s+imjPkd0LD9YZwjhgRJfElxjyZfEFzEIWjrsv/lWMnR82uOvPvCk
nRp5Gg+mDkGkEfybVyCIXzio971dEsQvTe0cBH71bc5oFrWSovYsJsN3fEwU8wFM
OdOs+6+9JC5MH7z5mqo/QLQlko8BaDtNh9uru7tF6/1rLsuXex2l14A0c+xS3CMw
468w6RxCzlajCdZA+kVMEo52mS6D6R/UM86lNiWIIDw2nJcBnXn29jhsmaLyrj7x
kkyLrVmfTgIGdeaNWtmr5wgY7o9OLJotXddTi/yqxftWFQawRKpjGlKVj/hhVED9
ToRCXRqdn2MKSPF8+EL3vx5ETnKWrbeVhFIlKNMx1z8jOAlfvXIBNs4neUpJZjtN
xz2d2jPJrCLozj7Gf2nWfqJZXplDHQIJ9C5EvaXdNMlkphbpWP+FIE0ON/xSq1M1
vUJpUe1p+/Nf77O2gNcKS3yTi419GhK3rLwkhYw8kqywf/hsM+0F/0nRJC/UgrSH
vn/gn5xpOXz6O9Dt4fGDYg==
`protect END_PROTECTED
