`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QF+fB7okFfFcEr0g0o59J7+yNu9LGLjSty9r+5Go/hiqwNOOXpmvonwl1DmnGPHs
TiCNstJVv3E7ta4f1A3NH+mxRmtudNWPLnNGnfk6YSW5o+Z1ewasOB1FgXgePF/c
cod/TA7pOKE9eiyfFXd0fw+moev58gNOVP2hvRstV9yE8t07pT/fO2ESAAiI9AEa
m9yxyPVI1dfnbALdGuBhvHlAyWy6n3vrFQBEVdrLKdZJxhvsSlxRfkcHvPknzGKB
AKu8C07vj/TlEXNpFXYf5b59OvxvilMMHvYp7ssfvD6oveJZ+Xs4qlRTXwkg9NYW
pShd0z+L5kDjdwyoSt3OuAMrVKJWvY6k64Tg/rz1XU5cgjh71S11nUSfLkqNmXoD
6Gk2d90q+Fs7H3mt9LVzthrCcV9/dQb1yec1+B1/qw4XLWRL33cYBrpsuIyCMyl1
Oj8ba+nlHRE25BDxCSd6wU5mvDTeVaSmV/5lOt90weyIlCyn5kYkUGK8zdeJcQ5V
KwiF1U67U+QSN6RBkikh3bofIGlk3PlqdIZf08T/R/kL0nf8IbxVojuFQdcCKkel
5Ds8EFlWWhIQOq1dv9uL1uJ5hU1tg8Rmk2cfLNL6HbqSAS8UCj5CnW5iRY1Le/Vg
KqgNR213sT+CjIvngHtuacaauo3X0pHrz3Sa39jlXHPNCaKVczvOvn3kUSPMXK6H
/AleVmOitmgM5y4yvXdYedAwyAoixu8VCOIML8QoaXUTXvWOdA7zq1CSe7Avljyg
0fQJmZDOvPsEcNTApxidmx016aMqrjhfcyWh+zzE9dwUxkmFRLMxcQcLYfBivgXN
9ZO9ZqH0ZHfqaZdb9GAHXuiOBRTOzryi5biShF+i8MJQgzVGeVounNgZOfVtHdMp
YEACizjzItJuluVBaEtY0QhLzkCViPuy4AQVfakjjMllBvxh8LOhv98ddqPqn1lZ
y7906VcYqMEkg8mGPHjbbj8TcxbfbwIwauLr8iWIa9DXNeQ5RFMUUrDSNW0x38cJ
ctFsMYAPq8FIO/jdmDAGcFWPNe2ZV5lI7Hk0foiF6QrciKvVVZpCN2dZxMxchmOR
RD5h/928/njTT6IBHDmwjSTGe4FC8w1PYr02Ggpws77NmtFjmNQXbrjOMQXWoCAI
CtOzq80GH530u6+8j7qGL8GUmccWCNRrewbnN05WW4lyfiaDspbP3vM9cNrv5yGv
0EP/Xr/Ft8ejs0eAoH/30ohwgvsJriD9VENKFFHThz7FufinEWPkVe8OVL0fGj9l
wBNgYCpQeecusXqqPhjOWeyWzt6lfAd+ZcpOWYQ0UQFSkiJzBtR/nVOU9OU2sXNx
xzX3zoY15CH58VjjN88m2Yw6HHb9ED/ygNiGnLRyhab82SkKxSoVm2Ih8UmOzp7g
G04T80L0H7kWpaARrRYvTa+jP/3sQOUxJtdgSB+vYfi3J/N5m57sd4/AVtzQv7Us
emmw+CoNozP6OCUihx2ScRSuOmDbO4zmMLsTgGdrXDNpTOJQ10BBUDSjfjfP+f69
SBYaCoDNtk+ZIyckLWz/fg9aLHETV2eCPxFso28H4uXGAAyEn3V2XvsZ1NaJCcxq
zedM/xwxtuZVdUav8n6OOFG27QajDLJZ9LyHY5Y0gpOPAc4U7yBa7QA1IE3AEN6Q
bePj9zwZ/XUxI9PB88rqMLRpIWe4r7mJIwmQBg7lfpQJA3QsyEo1u0tXNcuJx5RE
GAu7xLvIHGv/u+2j0mZaQtUKNiDRDANcQ+jc9M1kXo0mHccpQVnVDGe+8pkIpgQT
+OYsgEnkJw1omj+kaAs57+WWa4fM+GS93zZ85+neZVtlckV4Sc1LXJeijXhTKdR1
6LRo69G6uzi36ORr304rURtB+rA37duTjbXUqHwd2cBnqECYRoveCXGHIdWuAgkQ
yCFJPNt6xf9kCga5E/kWcLRRGg7KAlXDcQpIgN7osKo342XeoFR5+ptRv3um6I3D
wp9WBar72lzqv7SMejzRvTPdK4mFKHzWozOhc8bO2LZyu68o8EoHngpArOJVAYpL
ZJ4Veszt7hYlRzcWENGc1yY4tUlk6tkAPIW/IjJL4BdXpU7Z4oso7EB8p5k9eNiA
bumXImJpjIw69a7X1ddOvAPaWuFs7mZq8flRji3uvFx9I7m0nhzbwEYZ5o07C0Ip
3AkHejePq3RIonu3VDzsgppymI3UcM1SiKgtSWY79TMIiEL9Z8G/nxUSIRTQe5/R
3bpYkHa75f3cBugjOFKtOFj285rsYdlmBRb9Z+1oVQBVVbJdjdAQdgrSVGTTPRVp
EoyUnjvwrVSTiHD8vY2EJ7YhGqgoWPkjziop9Hn+cHkmnx1V1XPk/CftohDkm6lj
3ccPnvpmb4uKVR3zf72FVtgcDpSCNSmD9Qeyq4qk9DSfFqojC3zLpnZi6VEP/+uP
q5b3YDKEeVUiSDenaAFBSyfH/ONF0fwTpYh3hDU9xwuMMZfT2gQ2+SiciKUWTK1S
SFsxyQ3con8m6T2Xg46sPxWXFjwDwkBwbouNuxJ2klbwqre6U/UpwqicqqNFORGV
vLZlIBUFwptQ2wFxnpmKcaF+dq0XLULdoFaiVF49Zo7pEga6g1K5PQ4S8krg1cnt
z07kG9LGy1w0V0e3QWpfdjmJph7axbBWI/KtE7LHeQEvgystuik/S4T0Whw4fz/k
YRtQaFrl8yikH4obFKoJHeBcus8m926VUx3V4e7YIHJHemZiP2iZGu0G7XqyH2bS
rC2re8g+KS4sl3p22jVdMqGq22c7Ip5l+GtRS4J8KRPO1g5oKrn6IwsCj0NyDoQ2
S0F/LVL7Y9wf9Xkl1hx9JX1GQINZyDhC/5TggYao4oAgdjMwPHQ0xuc/6Fz42XWN
oK+hQZvKA1oGfBLJBNpYwNVxnYv84w9bunU/pMqEnUaC/b89Ysj3d8TnY7xIJcJ9
PWyfzday79UhS9DC34EHFLfU9eTtPozWgkEOM7Q5PyaJl3NUU2iXJfi9mPTX8DY3
M19P3NV8jXcaCCji800hH07IU/QeACSabnWWtRI0d34klKlhQqeml5XukjnaoWEb
siyA5huCzddfCtDI0SwTgR6SVWFoWb3xz1P5KW2Jmq2LoyX8XzxNw70OOSz4H8kz
JqcmJd9BbESOUJPf6OBouCJy84DTqJjL4h84UbYm2WsYDjahWQF+AsuS9NLPoWaH
9+Tp4h/v0Gfefx1jNghozrZRlKFQ1Sq6aNNDYYVK7BaL4aB/xnt1KCyRAQT9XAHh
wU2uLXIwwLwiSNc8CnbvKxGYKHi6lJFVhplHlFArGj/SQJjFS1bWH7Hh7Z+5DqoK
4AwUZB/3aEQMlMB6agG/nY5+JHUFZ+6xzgbuwCNnl+fXdN7RqD1H3RDxXK2ZhUDa
TNA3OKkSgMQrulyoMUhPE/l/Fon383PBhhQznsFo2zvyRR3EvqBL4vSGDTA7A8DQ
2RuSiYjoUpLNc9oLKgTmk+K7qn/4KzXu9ZsqIjD5yTwrIRXMzPY3oQKfFjKgOekn
ejg933NW/L/mn4+/mVKnh9xbPIDIo4kTK6IEE+9dNaIKDWWlAvXBMcAL40yM7F72
SRosp55YMOG/+MJCau4RDdYN3y9gDjnT52/GNhmFSEt3jM40E382EMx3hgxxngbW
H1sLfGdSceaILR/v6JDh7dw6GgAWdYsseuupoJg+Ytm1O18m3+raoZGpNPv6x/uC
NE+mpVWMSdyoBD++iC0dS5a1fXcMm/OL5dla29W2Zxc7lO6kgTvf0ZvZ872C6DgF
uG7YvaGQRQt70JjKfg7vsQXLONegydxEWHU3kCssIVjYJv+CY0ig5/qUCJcpfwAU
DtZpFHvTYvqfv3FE8K2dDqc60U7DwnNBXDbuFn/mYbfMqEoppIaN02qGsdLCFpQj
yYZhXN07+QSKs3IjAu8YMIuEzP3H5GnkutjWwef+NTn9tFyBKIsZd2800eh0HnUd
nlRBBLwPMkgv8TWSr5lNZd+gjg+djpH2sRmFCjyJCrInrKbBc+seYbWqHLHv8Q9F
tgOtovfwpsyHEkTuPqART3DK2w6AOZf1ZEVMB0ClkIIRhMuXjoizVGM/ggSqxsFC
nmq6Nilw6MpSC15KjeucwmMN9hVCaEQsLTnAfS0ofOKCUk6p3ChbRgaj+wQzhCz0
nygxO2Cj1HMWf8I7RSzt5M7TvepMh1/n7lCeuYYiZ3qbSfTZxwpKQTx1aJ9uq7dX
J3ov9zLr9G9dvZeEvdj4S7Zb1AUAOXSbWsN1O3/ZVAmtVtqB3OkJvSkvuy+rzP6n
YSSqmdQ0k85JuDFkB4cAETk9FJ2BmqeHAw6iM4C9I4or+KuEtklW3Cz1jrx3N2lX
wpvIz/SbeDK2WfLqbW/g8lWAbWUfypCloUH6Hg/fpq7mm/DWCvN7DQirPvRIVryi
t63puFZ1DF/xcOB3hmjSoVD3NOTtSQAm85vJd9hxg+xV+0YQ16scGyDPI21NuStJ
4O0uGmihbG3dcMaeABGKSsII/wgqrLVi71FeqIwmwXSsjhwoUld0w5YVRGXjJu8m
Wn3L9NHPtzJzX+hkRcqp9Ui3tPMtweTTGNbMjnuGjWhzexiKgQQ1C531QZj/bNF2
JantKjdxZlnMRXSmSPE7OeQC42V+k62Ud5rqVctdDHRqNZ7MQ7ZGNzFNiRXPb0P+
V1xA+PnOYy0q7MdHwfRjs5pRtpF5O/rUGExg/doCHZaJpXwDhXbTamaEeAseLN5w
0LMrUSkZmwMyT3PWDLm7W+iaCVRk6arBKip9UV6ZkVd6DAwRBsUb1TRY2UffCu3b
PqLsb+bu4lg+A/ll8zUc1qf9CqCbx27T0PFBFBmLN/QpOFMemZQ4daQUkMcVFesK
ZTHP+ivwJy1s+n6/D+a/fvMjFyBrm7ZM+lO+ADRb36nUv/doNQpsCu0QHHjCpQ/m
ROWQeqaS4Lg/a3YNinnGGGUWm3Q3au2W6/bda4tf7Tle58eNBVi8PofUK1lKpMTs
RGr/eeB4aIo0RUheptKvWzn7f/qbVwh0gUJpY5YP/3WqoKOCmMlLjfVW0UIZ8N/7
YChJDjexfBwkvnUd72hOVyhC89kL5t+5KxMx8XMYqaI6s6CgHk56buSzCA2uErog
w3fvMrgsP0QhQZyKIA164mANo5nqPqP+lNb2uxOSBJ8ESQuO4XRTtMOezjvNiG5+
XbAJIOgvsqX3jVZJaZHZ81yAaEKBbJcd5k4Mimx3FzpBJYr2fqqFpMH5IQO2LzgJ
OC1PPfB7wh4+s2w/bW41ehRWZ9UV0C+xo/iAKxs8so4Ptk2lNGv1oCXD4k9gH42R
F/y2Z1lM9//jHpNjPYoMQuw2kM2CEsGV4uGpfsPyNo14oN1zf86pY4y4OE72Es1n
NiRzz/IzsjZW3NYc1RlxeIkCBU0hK6mh1s4LpS0JMjgEevQRS09X2A7Q5URxKRFT
N13920OpnJfGluI+r2mWvGT8EgUsCT7Cnz2MSHpBemPPFN5nOk+FglquIO+VQ28r
ilh7uRv9wK2ZF1b1fiN2cV6H9xBl+b/jp3uECFndhlJ5YA31RWWDpdHfOBZi7UQV
WBgxbswmZMgm7g0jFYYy2FqUoi8X2Yhf569NlZLAKKwbwKXM2lLzkO4PocleVrG2
5G2GbNsVw2/5hxB2pE+M8JQ77lyH67JD+mes2YDC+udOtUR48qtC4jZrFNVWu/If
R/rw67fmvstlmAodeepclGj07BEe6IIlsv2ufRpPdar5Luw51j85bZ1YEYvMv3j9
hjOD77rDwF36FVos6hkMnv43m1qgz3mH9tQU4TsEcJ09JBuXKKPcENXsTt3PeDmS
3fxwGaHEmw1ppg7rUCE3MUiUse52vZd95BQ3FFfewLxSEnjX1mnrW17B3+HC5Jrl
mqnbF0IKyJW1sSOLC6WgEY/TR3FP9T4tyUkziusjGl4cvS0hbq2s7t0qyXkDN0U3
qkSHZw++H+M7TVqPWU2IGN88eDrxvlvaFCJ38c0If30hG0MVv17r2X2nhb7ICA+J
iKpydLsppVt3ybPxHQVYvxdN19aGRjLd8AQkMdMaHDs=
`protect END_PROTECTED
