`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HSfAiTqnjex+eR0S3+lW/sBz53kkguOrvdgdIJ7p4iGPoP1Jx3bPLpSU0fjg2kQw
2+gT2naAxCk8Kgd6ZyOGrTR973HT4cOw7y/7E1J9PG0Uf/odYi568llvjBw2Hbpn
FwxXcLoFYsxNCstPV5Xt8LHabXM3RK0v4dPjV/VgQNkFWv1Vk1TQ7BC9h9mF8CN/
UPSO12xVzmb0YOwTtOxIm3rM4dXniGyNj5i7dQXhLsDNQL43T5twAXN+R5R+RrM1
YkIn4rwX4iM0edExZgVQ/+rFieJs7z3d2EopkggZA6KEOBvLclCMDCjUKlae+QM8
GVzfEHAi4kFXkt+8N4Wpr/gndGJ3FU/TB6hFZFSJFSHAdMR0i9mLOevM06T4ndmL
D0j1gMpKOrtZuRWV9BZg5Si1ujNw5fhLLgT9j5cfNr/COPPa+FMj5tUYYeyF4/in
zxS2u463oqCQhHWYALWDEWnHsPL6vGZ75nzQ19uwMruFWM80H6RJciyKiAWLouoh
Bee7F3CcQNF/i48+bfOtW7YC+EsuGZUpA0rZWUSHd0CN7i6iQZoHv8WkAYmFNXHJ
aPN+iAeMz2/MIcIidJsYUJ5t+fJcUWPGn41gACzTKELE0L//xyyGh7WEvL5pYObM
4rd+/hSzCz4LtIMsINP4BoQ7lTJy9R1Ll7SA1WgbmUxHp6qJWVeXBUHnOdMx5CJN
AYnqjn0arKXg0Wmca4Exxsu55sQxD5WGQJgv5QCE+bLGjZyQPUQIndqQKxG15Fks
KbyRjTGsKt0583LvdkO6PKTS/UXGMVs2QU/llhRQ4MEujdgOY/LIab6zDsmcsnZy
S5H7P8OHr53/YNvOnG8MIr+mLdz9TQEtWRdIb4rvdQ1QnHGJqf876Uluvaxx8RIg
AzyexjH103Z6RiLW9GGu0+reDHOf1G4Wn0EUjvfU7Xej/4+o44zEXzvlro4iRtg8
3KHHdq1Q8dnnjv6kEqjbBGoHAuHBtFOG9rPCDpgZYygivDPmSY7aokeuLNbOWkDV
Ld37P+HC2PbwCKgJoNyHKqN507l/4XB3bvqR/t7iCt6mxkijP1PIJvcxR+ncgV+y
Mvyp4mJ9u2GsJ5uIMCOzdIf5opf9fjWe13I2WV95fj3V1W5rdwOcp6ZrSsG6IA1S
RWxgrwnYsTuj9hs25e+CEJIFD3cPX2xlEZ/jtczeJxisLdWNruHN9ml+TZOd/Iud
Lq3ytKYsNiCjy43izeOpAwXwLhzhIBJbweUTAcA5n+gSFVbfQatt7vCEhcZXd3lK
z32yMTGHfcWfTfIFYFAXqsq9Sp0fSHf/Lc36ewvj6dPIZwGf4r8uO0IuE3f0vk1A
SAvsSyz5a/HpaWbzsluHYkNj9oSV/gSWy/I5gxynJqs2gfGJle7rtpOHMku3R21b
2ytVJi5bI3MZbH0loqM5LwJqmXXzIXs+aCtSzbnvxKRWnnT0dezI94YGrba/qFHP
Y6iUkACWcsYWhBSd/v/teLYtmuQJ4cA9CGYbD2FG+cqKIXQTEhfzoDHFIqq41Opa
wNW75yjqNFFbNJ30NI3ilA/lUKUHp3Zc6b7HDXALDFronsAlCyrf7BPXLeTcoQza
a3mCs6tU9uLmCzGQXhm/iehlneROrr9wKIyBtgT3BBZPRoG7guYqaG6KUo6fZQHv
Esx9heCcgUa3bcIuYJj910qfoTQHp2Ykt2d4DGQYgMsqhOGyc4jLCtospzuEgz9x
9Uxzu6a2CvTJMXllLPCy2fU241pfn+SF/Ra8DO0ZNgSxExxzzI8EykzMj4pptA84
r1xRbeOIFeH7FIP2uERahCVeAk4KO7CF0CAyG5bhzvIUiF4GeiARPoI7i0krXTcH
XuDHxyuFQZZMmZOIxrYAakHd2Pr/pTsPm1aCJM8OWW6nVnltNdofNVB2GPl3B633
k8s4tGHjEIZ7Di5fmNNH+xo1aNIh8KKA1QQDtGggxuzkm7Lt7aI0f+dHfLIOj1CL
j+/7ybf9r0bPmvEC4+vq1Avu9z3J750HMeQsT5PiTem4JrhG9Gf3t9hfSnBradzH
NhHXl84E8EqKAM0kjm9BAECkpqM6Ty5LlbSm5pb/AEcplxVsdht4gPorpaGf/zIx
sdB+yKTRGRWeSMtsDf7YQoGsYmAazzwp/caDFnL92ykJ/Dp7KgYysywsvg+rpKfz
B8UHF6SAMHwkwdjVdI2/vE0Xie/1UASJChOKL2EJ8rRBn+oLm54TDXO7VVaSgev5
4uq0PnR7Pa9WOurqc8Eqr5WvPlQvc58GxHZvWhxhn5uFZIu41E77bvBHjlzw5jI4
YLsYKmOILyYUi7noJeos4PcjowKJKrWmo4YE931qXotBu0mJ8I+DNk6E+8+UVbqR
/I8OC2cH6PNhiW5mamVaBssfcs2ceWdxcAW3q9lJc84STEOTkL5q47FceZTcNv6R
Yy4QipxK79y6cV1CXa5K9lXirgPGlrie/abJ0Q+v0vNb/HoEpIdv0JOB6zXMkoRB
ivnMPgPzvPOeuYPSL3TBxBYzTtW7Ymnx6EMhWpZDKxbz/7bFDzImsflGpp84tz5X
DDx0lV42TVJsLPxIY+8Vr07JKwnSYUaux0Xa+dBKv22EFG4TGsnoiHNAjGv4dNWR
tktrszRaoEYvwlLx17+mycWkf8+9LfA2G1spUtdTIrjkVh/Ph9Tyw4uo+eIvEXG4
bT97+6A8F4rUV60o96bWGbRL5v0rDOYssPniQt+HFD1NcbgFGFkDq9t+sPsANDcR
5tYNNlRnBTqMeF9NWzeE1A7chOnZNJrrMmENwDIhBPF/a/L+JF0+QY7zBARkM4yT
QooUGuBd9ZvosB32VjNuHq6t17coug1RsDCEohuGijFhoiV8rm+OgyVYSWMjA/Qa
UxFmd8KnmYMpbJbrbf8EEfE2ea9lTjxfsFCKzZpNeG3Tkn5tYvCTUbtVotSNyKTq
prw/kktxn3nzQ7GJmWgXfP8Tngcsr1t1YxFYpC7lPXa/CBDUfG4WTXzB16G1EqhR
CI4AEXKch5aTuQ2eJLG5+fN4LukrJBxzy5s170QdWBnss632macYjpYYeNrScEDh
nb0SJDBwPx0PFVHJZG09xEsIVnh38NjFP7lpEJuwB65xhY6Vi2ajqjEy9XTiiTnh
X/wG3OZ9DqHB71NsLQ2nGlk5mOrqGeckqOyFz1i92OBq808oQOn0vbB15cx5Pq1X
A9Ub6g+Z8+BKsi/zK2cAGFf3aei3wqcncRYFIPbw8ReGR7UB1nGIaUaspWwLGEzt
ikuQfNdyiFMNRaRxhjAUmoVgedXy+4Nf+bcB7ScsIeEPZOQB+CEbZ8fJGxL2Sjgf
koulwhiFC/vSqukYNZgM0fJRb76k9Z6pwttZIVCCJBzCKEZCK/CEdXp1VOifCMUv
EZ36hyiOXpb8DwnltE5l5euibZf28RUCkqxaO/vEw6I867rNnMwtu7fqqTqO+LUz
Q6Ie+7Nvka0R4kRUVk9hCnf+P1yXVKyihSlVB47eV+a7ZSeqpEbudk31aHNVdSog
WTWEVxmjFCx+KyJt7sPAc6J1V96VxW0xfgHeFSjh8WpCCELXW3TQ/GZDn4P+Rf7v
dBe6UoyM3oQYH6jxsqan5t6SVyhyDvM3rSf42fvzkZeFnQleRpHlAMBPJhaYIHjR
WuuKjS6URiJ2YpXwNFiXdjyP5wj4Aw7R6wdW6lSkvXtx5dLB9S3ky35vG/ZevkS4
Oxj51UQrfmFZqZbEvqLmMyEEOSSZF/ZiCsbqRE5aKo8NigQufcQ6Hp7c+/AkHiAz
rDYnrPsrAHzG1Xwda/R9U5EEKi8S7Ta7MztUkYVVkgaM74E0uqUWvd9jnPV4RWdr
XO4dtUHWtvDJUb3w6toGNqcenmDv4wbMAnOTQPDTLof++QXwP37rdOFcIU5NxNz0
lI68oR/8OJIGPDyXxYrXExHt4hgnoo6tKb+bwJ6jJ/4RhM8ODDO1YJZgfVUAOp4U
FGMficq3J6w2XxW845ZcYld9LPAyoULZk8dG79igCxlki3X1dhEoh8Z1LoCy/V3P
Ru217yBpOku4y3Pj3wfsbpSIhIz05rrOMTXwqYlFxjEj4XHCzq3eQH3WO8i5zZxi
C5ziRakT4cZXkso6Gf7wbZwTYgaBXUz/nJSk/o7aHrLpg136IF7/Xb4qp1ju9dhp
K/Zk/z8fLbJHiL/lnpLSdpJix2jWjEXeL7bmuCsjPBdXLedPv/HHnW7TiwjuyyLR
2S68A5DALfZ9HY0haEQwZ5fPVBaJ+PCRLkBs/o+ab9iWTyJ1SX/jrxKWmNNGat6l
n8G5ATxOI8Ogi9pIK7uEi8WOyTQNoeTytgHwmP4BBhLqB7r1oEOqwoAsruxr9PWS
rg9kZquTEPEpv7qhBu9+twZzujuzbzlR+Q0QornaDQV3ldfqWZKTtkEOkUuHYctz
0jjH+VGDZN+Hsal5qlrWabc2LhkGqOX+Z8HMtvoqDkS3xRoR2BtHY1YwWW1xmsEO
ztG/+z9AgU9Bu6b6AatlxIQXYTHwtg1KKlV7HzArRfOeH7zQqUjXGtT0TkZaD0a6
IV5XxgL8idEsY2FoYsgjzDoYYf8vvx3kDLRWbWvP7c2BbCdRLXHTSnu0ioiKTVIs
A9VLWgHfaoxiDjYF5vKogKotHG2cRpgpNCKBKEHXkJeIu9HbNCFmiO/G8nFzCd1p
QtfClcdw0Ax84T2teQUWMr9Ysc7lcZyGitFW9VPWvbVNxrMuO5DowuNrfVYGoc69
NDVCz+I/rDrMnKJkZINiC0I9nHSD26gkiqqkWAwQYfnyuVzwBnPZLKKBtyDJUTe/
qLINwNhUOpw2udei2DTKYbko6k+ghyZbgfnW9lKmxHQjulcJy/SVYVFUzPU9HN9M
LtYSCHkXmKmN0ugR63j83ioJ41pAu6pK5+qQi+2x5gLWi69Tg82NO+2eVOO/15iU
oQ9CenTZ5WKKIZHdbGabTzJl+8aJWP3ZgiImastNgny8hfBtfP0q9eeKoaNLAIcy
mQQHlo87G4kriFCvCBJLCWGxRW5MoZzmEGjCHpGvpgb2cYMoWpvztK+z4zLZi14g
i0cr8y7eFuKxZBFXn9yEONXuKV6K0BtM2BoTOu+nI3snjjyy7F+mqKpDKgjqotVM
B847n6ZBqbEcjxsCXPoOEHDt/HMUUyzdD8cNYF1Ue7pVfH8z7tbvwZNalYHkVijF
A1AP9Zric8ClDeeJJn1elTwAgpBzM3ATV8h9SChTgefypAHkMsK6MRntZDp6SFnf
bzytMtHbRC6+AHh32GNTPnpJtu83yBZVzxQvuv9REbLCeyY18Ujo047uxVNvbz8V
CNR1LFgj3u1UUBsHizuhEHlPfb6W2mIRsN/SpDiB7KncNdQ5kIUQFmcCFP4QnwPd
88ouFYGNzPG97BsmxB0QALLlO9HZxZEP69TjpAcpsU+bVTuW6jVhQ2MRsLRwF/Dk
uKc/S09aEvxeZiXMdfkf+aii+bCqFClaC2Z8cYmPAbFcaNk5hvpF5CKiwxoyJIoB
2TxSNUA0qXrvT+1fTwMkNzAJ1MBMmwg7XIiYtblwQ+56hW0qM6nQvE8Po6vxsdHX
bYgS+i1yDNPpPrmC4Pg+DyaMLDJf8FeFvOgOK0OjFymCCBrQKba3DoQqMQ9q95mr
eflL/K4Kbg2n+30+8Hpjg/xTp3WcJoHBIoC8QmboQbbliz/3VuFelWuPxJRk0ZO0
TdoZxlEk81TfSG0GnIDiNjWv/dqCa+HOHo3U6AKI8BKN/0N3YsMu1AYWGYIKWhe2
hovZe8/jkRABuSxf5NA7oipZD7MNyYuAt0hYvINpwQ9SWHT6nKS++wMksxVi3j9l
ydI2wSDp4UfB0+EqnT2OH7S7efDt+Bky7kBFzW+DO8Jo/P3yhAkraFKMlhznsFwb
EZhApR79euSXihWhQkrvUawqYogGhQNfgrfE4BAuE5f3jBGml0PJ6gbEUWPWO+pb
lfm15DZsjPl7700ETqgjgmmHKclVY3v7V56rEkWojRWrXwLLQoTX2ozF+TTytPC0
aD14EMbOYaV7/vNKeZvIFgBAOnRw4jbTPs48XP7nXlY=
`protect END_PROTECTED
