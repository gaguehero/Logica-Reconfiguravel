`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1iyzr9WAG2IKLVV3P9YQ8NbhYotfgP8lJ2G4FRlzU06SgGGEVn5l+PFs9r6F473
kD3aFrNVvL9RtgdR3kBnh8fbKmKcy8QuiGZYZiAqMlNl3dLsU1H0kDkxHvkC7nr4
p836T28+MFg/Gkjs0qXBL+PVoeVNg7IZksOOpgykYQMc1TD8t3i5+zg7R7fo9q+d
jOV7ZApirlwcFoRnFk3lUE4YSUxOjt4vdq3SSG1F+5AA2s2qpv5hiudhcYEu3Mmu
5x5Y3CbKmRmH/Dh0CDweaR8RBRRgxHchSkHa6qdPKLZOgWzXmG1PWifPvBY+CHsg
JK5moJwmSjvOvm37xDAHtiDcZfNkFARt1SwqUWp3+F1dLiq74ONjpCIPuqxPVTKy
fq1/Lv+LcSxkPWKF8SJpsNf/fVD3/9txCMUb5xPG7ZwGw0Ju3HkFD+dVOms+cmU1
yEmQXq4cRh1hbTLzGB1Kqk7MLO2jdr81c4M3X/9qW750VdeXFtQcUSdDNm1LSGcq
zIeZ6Zv/jao0DMu0h2k4UkSaAwhQ+123GK+JebFIbPTxTsGkCr5DukPhXgIykT6+
+/jgpRfE0Is6BAuQ1HePNxeKWJoxVxGBaSY7SykTExGeFuDD8mmsym4oY7Tgx148
YiM69fx+b40zFkD9So+vBugsvGwF02g0OCJrBFn5y95eRYOVl3vM1o9Udgzq5Kc8
2bUHO6PBBM12XTJdTJ7zWYVa9ysY9MOSnWtLcKlvmAtDjLoAkgvRUMvngfMOdmjf
WUT1sOTAl6kLQlvv7Sy4M21UVa/ZdezK5jkc+6upouaDSDeKeq8S2KY01q2JQfor
BDKytK57+rrhw3Y1Wa+9NYsj4+udv5WG4Ym5BmfcXDSQb8xOhgJPJd3a8FNIGyJy
+oYh9XSO5MbJ7vSDBfiqAdo7W2H0E/MlHkS1V/pdxJgBk7FPHejWzPUZ0yk4gW8I
QzYGqXAU9Z7gtG3Py+pacuEp91x8S4ybCjiW6sYCUGUyogGVWUeWCgoydf7dioRs
WwCFfspul0+dbU7oMjq0S3oayS24FxCYkQz6LvQymPzEP/HNecernRTs5F4+yB5O
a8FUq6FKbRtNslQbmu14cpZYyatoF2dn5RKjvLIUTC94m5Ep2AB1CbWMfqEbscZ0
H9jI9HPQavsqaHa51ZgwZC0v/3xauii+x7HpBCFElTSMtcXeBBBsnwdHV1S9nv38
whSnNI/UksjE71mPJyKe+OTLkwdHrK7DseB/C+PTLRBvX7wl9cSdJDDJhT8GUuLU
qwqEFeE4eCyfpPrpa4RbrVCBFFjKnJDKmwPBnCDffWmCk564T8e9jKfzGtYhvZ7p
mvA7Aez0d1xJ/KauYg3x6msvPpaTb5hoOKq/pawNOwyx3fz0zFh6WllZzP1wsYpa
PVUoxB9Ke5479yVNOlZ0Eq1foRCVjt96Z/koixcy8JDHzaj5OrqOeXwxaKCjb1RB
hQ+GA4tT9CNBlx5MdMJdnZYtz9Gm+IGIDIkGR9UJFSum4/hijwAeaEakWR/PXBRv
dzW/l109J2KjvJQzgK6WtLqMMf9h3BYWq5spZdYg1KuFsd9K3SV2Ev4L2TMjLIAd
B35jGQLOJQe9wTzh7SbGK5kaJNFYN6XaVzCvOB6ZfkRWrVAS6gM247L3lJfFhmuA
EST5e/fq4yApsOifOmV1NKT2t2GHg+/uCdsY2Q2Z8b2pFj1UzeNv5jxbImrqjmQM
66HmeSogIRaEe3rwQCHhO3MtH0xUViaGv1/iBHwYWlu3Ms6uHcQZK/kDWaDOHnYh
NT2zK2kGdR5Bw+HpouHd5rZAXtFtfTP2obs8DZq54FPADIT9FMJpUgopiaz1pKI9
Dpve/eXjRtakevLRalMcx0bWxCD7JnwFCIKB+JWP+gsuFYhbkk8X4ISoDfAO6X4V
CWW9SaYFZMRvDozxszJKH667SinglPGFUgCYCffHt3Ew9tnuHr8ewccLfobaMSLM
PzgTSD9ZaZdU2Q8OqcYpNcpYI31wCQQwDMbfLj27q8r2ltX/eZYjwQuTqVYLcIO9
tFbIUCMvcWIaEv7id76rsgCPt/k4+toMRzMFFpRhcYmUIrCSLsspS+Ge8DYyrrNy
DQJbVNRujPwSvgwOQvGU0s3NtofeVkszYJy3Otcbb76Jzk3n+TQcoCmShQOg8ivd
Hq0kK+gL9sUnBJ3pVGTvoVYhhWKdlQI2Hk1CntCRzS+hBxijOZ4q9Sjo7cuFBUUu
BSFnsIDxdJnKTXBHzsvPqQ==
`protect END_PROTECTED
