`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hpf9a+wcNBqXCruLIO2zIwUf7YZFKHl04eKHelpGMao4Cxxbi2FS1SbgBg800RmO
M//5DveU7ZwbWbJQ3w+FJiNr3DTrytDjSJgNvCMpoKhPVHFPSQ6NwXUJP6OaYLI3
4nEBzDUZgbpOzJLiQ8s1AMKQL5Jzn9aQL8liLEbP0jVRrbcDLeW2YAxyj7Ij50DB
l8/S7qufpXgnVOQd63Nk00M56y4CxkkcIuHWl/KmbCMXWDSaQoFFJP514pTUGF/r
eJdxRwA4Pkndyrjo9GIsAKXiAASeWGvMJJaoR9e0zHRzeKuJQL68X89tnA7oyuq/
flBI0dpB9ZQX8dtcIH0OVpzSW8zqoIuQj51whC8bxTbVVJxXnqxqPv5AyOHaQZqb
m1+onfJaNG+DBOR8tBs6u8M2Swh+aMY1B/zgNd6Tm7r/ufnkYKH1Xx1w+IYuhvlA
ewe/n9DZeoitbWpQqyHf/7jgGgz0FGGEDUB9SZ6jaqt3FUNP4YmTLSFK0efWAFEa
HuzHTJUMs2HvcLFVGEN9KB44eK6t2mhS2Gls6nGGaByG9ptIGdFAWzwmMccD5Okj
Fw/XYUP2K+wOKYX7P4Xk9+xx9hkHVe1nLSNnvfb3/vOJiFnMpjTC75g14T/vBCgZ
K98D01TIzTn0pkkhLcIg/etDJyt7vBIzFCp0CNlM7jMzK6Z3Zfe4PAl2V0tsPS+p
qmTGExQK6r6TsG9Bj++YwNlXe7PJ3botWkCcgZ+uOT3a3rDUEbUsOMvqcBzKQhzm
4Oad1OtaBO+GSA+o4d2O8IiaGv1bodQjYdbPxq7R3mupzv9uQyM/orIFuUDe3m1E
sXKj67Nb9chv0AeK+ImGKuKm/WofdbRP+/n3TeNlF/xVVO+mV0xZznwGt7JNZaGt
Tg/XM+3vkh0mOIfDnq+ASbPNxDh6NzLzas1Bt4XOzlI9EMPDsvVscKLSBa4zJkwn
Q0TZ6pVQpjUIbbCbIeTnHZygsp+MuwvJBx7kpnDbcTg31iEMmGNJw8FqB0nz1O2a
aPB1EmvPwNjANOH4q2T6tWgvm0ryYgGJc+bEi1MLcMXIwRAgzcmUOgdbFYhZeEkS
nuVP0FMbNMsgv7QPa0yEYx+iZ0LndV7bwvFBHs3qo1+Fg9WGvO1L5GGPG/KBJshQ
Crx21WKGkCXcn+5r16T89Z1ZIE0//2xl5L52e3UDmQtmrnag2WWLVgw187LWH+U9
PUbKx1xXVpc95pe0nw9EGRHl5ZrG9VLtWQdx42ishpfKD3+s/3EsL9zeV6L4NXiQ
+ga8cG3cZk4fAkcwSttFWuD+QR8WqhEQskrLohXwbm351pVv5wEwqINXATHXxUMH
vsyghMp1PV9kWUnnqAhhh4ZTTUkycaBLcL9jisrwVfoPYGc1mj5+JupvLWxBqXBg
bHRT6/KTcjsmzpkZyHyTJHz1vcsHLFc6srnjVTY2GCSDYYgOhU3Q2DVeZS/Cz5H4
JewXDmenkxpbHH5B8Ezc8FgPg4yv/5bPn1jOtVtbzbXh7nCe1mouuqq+c18u0RY8
HdZw1XDbCIHydhCALJw57R6gpgtHNT6l7idBUydfTLsGYERil9KMtRxcUASjZKfx
8auKhbxaDfSRGLxa+LqKNxHn+m2+L1fBaW4V2DUxBfkOPxEa6lvfmL1EqYLH1a66
J/fFwC/yoDxaXwxXpNs0WgPQQyEECEhwAGWdA89eK7iRS/CichImtX67VpMz1Ziu
OXgXPh0CjKt16Unpy1E8NgMnLPTR2DyzJydR9VtJw5uL78GjnnJvm8DfKQnSSnYK
NM8qv4Opa/cic3NE2WRn5eRFSFwXAvrrjv3wSnXHRFxfogkjY1G+MNvBs7eZJE1K
6+M1rhqgjqYHh4ZYLn3I2mkTNwi6t00myeLz7d+7DcE8huGLfEkiJvSFwrKgT19Z
A08YnHuGfm2BehoZVxA98oeU/mO6X800Ci+FTUyyh+hk4xftdpUSc1YaSdxkC84F
JFCC0fx55wcylVj4/IDr5Q8fbcPcdFRifrhMP2Oj8iv2jk7+it2UPdtKuI85FZnK
wAXCEdIluF85K8fUbpQudCBLC+/eKoVSUJ22Ga4ZEVO/F1EIHL0DqLlYuyceUxJL
kKqDdozZ5rsUgUNixo3FTJfFEauJR+uYy57pKVZjnNTzQpweWOecnY+klnASmmdV
8U6b9mD5Dg1/rn8VwEKrAT99fnOtExdoRhxu7LXbWrryRLwnNiBUZE1XR+6GJp3M
M6Io9B7pJRZzMk5scoCiww==
`protect END_PROTECTED
