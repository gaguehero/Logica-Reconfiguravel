`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYNubH8aw5kZ2+ewJbJVq76tliIhRc4K4eg9Boip3Hs0H2UNviSWMbbvD7zO9Akc
KfnCdaFJoxEh8sR57lAMqB/q9LQkoIUqoT9PScZNtYpyANjxDyA6rrbPEcI9qS6b
YMbFaslqwELBejt4UB6hMQ3L5Xeeqvd59v4J22aXt4BiQJPLo1RFFzgi16azR72O
/mkPf3SU5rFoXBG2XtKLDg6fqobftVLddvuDljZfoqWjHWqCFl9dRPmViVonJvUR
TrwIDONxNbaLCSsR/xpp3/+EcJDoPrXK2F0Dhf5yeMa/txI0e1yjq/tMoB5MHwRf
r+QfEWgcg4Aj2fHVI6xc712rhENSCr/Ds4Yzv5bj5E3g+6KDFvmAMQ5G5c2dpiI2
P1S2GNx5BYPTlAh5rgos+3wyOhKUYbYcK+EaQZsY6ibD+pw99S1H6PgioejN82IJ
0h9+eBObZK+BCtj4Kpisc2oMQOzR3BeNSeNF/lWLhTJe22n9hDuIDEmHtS+m7LAD
fhsWPUzJisxjpR/TmZ3r6CYeOTbcHZhMtKuPSuB/ge7zD80JNe76DoxqD+cLmK4g
eLJnVUVXVatW2a4GPwcBPUjY81VN4gV1np6nblZ6GM5xys9B2vlgoPdNeDxi2mNk
K6PJFYsqqc0SaT1uqMI2OJ2BE9TUgURtMq8TJsYosh/eZ1WnUuagCQgfh8U70XTN
SPTQNrEr2cDgQAXcCuL2SfLLc4KEzrwCNKPoxqIDh+YYnfqItA9B+N5w5Ylqafez
TYsZ8DaMecuFm4ymVti/IEqKZ+7+5nEDdPYzTJnHmZcEBLgLQsX7TBiqkZ+3+cOE
7cCGrPzFMqszaGkDQt8rq3gKbkKDWrBGla/pv2BVvulDNLVVqUw7Eoea+TMpSAJH
VKrNO4SGNHHXsDsGjY20mpJ0/+6vHEH1G0vlWkGwlhrQUNc0ysr/SF0uRk0b5E7n
On9g5W/uxZk2+pKyI3Bwl4dP9w09ByKL/to9jm2DiDnLjH/wguepgPcrBFG7tWOZ
gC+7U142H6RBFgtbJo0PYmLET+n09wyjZBsUsfJhhETaTkazSAAyab2Jh2YGnSQW
ViKEjJ0EXH+mSxHJpBjLV/s2x3BL/JupSTdoIE32BtGHmlv1l/mxNK1Uvi+aaQFk
kzkHvpHc0y8RodsMLwKMQoj8JU9vtINKEQ3roU646bESzJkRwFzjLzGSRsSl8d7L
mOZQzT3pacIk1XD0fxam95/VMydvg/2x/3HlBZbQcrZfaMG84gh0a04nOdALeVGn
Li6ZclrC1Ql8XisrMjXI+IaHTIlxyFOv0LVwmII3at5VB6yMNTGDu1744nxj/Z4k
+JJqHC7YIn8P2tm9bRMPz1dAk3XheRZibP4rFGdWbfvSyirQvM2BmsWdo8S+FnDb
TT3h2LMEB8oBxh8ib23HJEJ5FgEPmW36EGTgSyQM6IB4sdLc57p/ZJ8j1r9VWnpG
OokKRjS/X/iMc1umuw0HtmSVuntwTu8szgl/vGnYlOREaFAyIxQrU2wcD2TLS5Zi
zsQYoUcN+1+sXIcpEOumVD28NpKVAruQKuB26ZB4xrnssf8pkGZXNXmcshaBhgiw
XK++QB8Fynk29DNKK1mof80K/hvtS0iX2y1a4pfVlcqwSjkgGJ3ZSN17VV6jzY72
FgjlVw1Jse7SZ+jdZovNkA7eKyoQ0u9jYkSIXzINE9JnRE65xT+WcJQb+YKQ1a5b
GhcmCeCoJfI/SN5RGclBxqffP5G9EmOk1J7v3DTpc1dev5lubF8eO3wDyRT0jcF3
9h+K29PmPoN2xeLAN+1AiffMM+2eDf4UWdYm+VCW3rPGkBR0MrmA1aBPS/ygSt6G
pmHdQO94TCMTmMHFApRnhBZJbqiSib/Dcn1RolLXglwTEOzO4iykJG/Q031FBLkb
d75kJgOExazAseY+iD+FamjLhyEsY/yLEIv+qFGIgSOhtr8EQEAKvIXkZKIe6U4B
mTlLff5IN01JIQ79JT0F/A==
`protect END_PROTECTED
