`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHqFlg6yES4Bps0fC6x8kM3yEXQYZGpbfq282rFF9RkcnMVLF8cs70vkKpQFFG+w
yug5AonwOgn4r7TflPN4AwfAWNJz3smKUhk7TvIVCqI/GXv6VPoU0zmxW7LwI4EI
SwBTr5sxYcD/Sf+T4aV8pmSHMyCXj5W/jieyl4Yz2ozAFjoIyqGfXXl/s6Bj3Chj
aOtKs6A/zLSp+EMZZhYmcQZTAw40AGZZLozwy4d/s8IO/4ns1QyTDq1TrmX/ki0N
cy5T/HRQNQ9dcc4JstlkpB35jCEMKiAmjEAz5h3a+9PfJCRqEJafihw7DLLhNclc
cYFnp25x5YSrrFETL5Qa0WjYJSsXQs5CySyKcRRp3z46HXMGHCl5Zjkd+YBsbDto
kB5mC0ik9FZCQP4F93skeRhQzIY7MMpkzOubegfuWkdH4xxPxM5z8CFbHSiGQmlk
SP3imcKR2QA9JH5cUBCMya4IkWbxI5vu0hRB9dKBiWIwLD/zAwCRgY9yMtCD20PC
TjK0dk56ZX4pn57M0oXblVtlGNXQLGT1fLZ/mEAVs9FEm9KQ3O9+bgWR4YpoP/Ni
HBE2gFVSYtc7b5+404rxOC5pZdoF0Hd9SJU3MhzGLseABWhOWmXLqqA90qwwW8I1
fkN5L49s6tJ5b2BSoXdp1BdLameElSe2N4su0eKnVnS5l1eF1m2+oICMToZ+4HXk
f5g8i18yrEWToBzypx09z1fKZUy4pJstXwcx7pd9xDAbWKo5KaSOjsRlQzXw9kt0
+1UsA9t6MbdwXZTTLAvcP8bkw7g3FDozwwtPvMQzvEiSLnQfSKwJix6VyflVwFMX
6oymt63tY9x+w3cJ/pbnRdTJzTqQ6vFnrJb6IiLkNrUeX2Co+mU3wukVVIyLeJi6
oAIGUEVY+QIFrshSg0euHHMm5PES5tVMDEVn54cdJkYlEEAgezMG5+mOXTQTNLRC
mtzp3q5O5NZzCpY5d7n2x4kbkqoQ4+Ju082fu1nwKuAtQfWNwHgLTMJRi62opdVE
hf3Ynpt1JC4c3e8lNi1OIm214qzyTPuSbdkQ1d9Kc50JZpC7M5CqfhIavay3uWir
ypPE4TV4TXRwwKQ+4sON4U1rtRY2BzF4vqXwnMufQU2wlesNiMeXjlQmgylKuS/k
MiFJrovjc4n3NUeNC+usHlx473DWMIc3sGfkaHAFDuYBw7TZvCXWOorN7itysD0k
2QSirG33bSUHH2dd+WyCQ9KZTlox+400DPmNoQZJ/dOVuW1HukjMJU81zOxKcXUt
bByO1Ui2YUlvano6ySdB2w6mw7KrAtTz17PRnY9Z0QjAZAK9ZwDseXFAw6iX9aHF
xEiSSDNyFqhof8+jHXJ4VJOG3tIFrNRBWZTH5EZXqzlcSF/P6wyShnKiO0q6ZQli
ftn3mZQ0MsQ9qKczz3FK+WCNTX7Jk0tJI22dr2AumomroRmbvObecHa1F903emZg
8LvAdIr/gJENIvKkwCirhDhdcJzqN2x7qj2soIEGFkVmy5yItZavQa+2tw4naWzw
Kt+IMoxzO/YAU5N2KD+NhnOcGL6ZJ9gn2bvEjeTyaOa5wjAbYvcq+maUwfiV0QRr
CGOy5C5UyGdGFoT1iRD/gqUgwCVbm7CKypKeJDHkBwlGAgPDovG5/lDj30fAsAJ8
zOmKL/PNNLdWUYt20M+aCijpBKIdtrm2Yys4rh6u4eB9mTWmfh5IpWqXVwQp8NzA
rvJe4duuqFSmUibguFMbeyazQJGQFiPr9HIYInh1eOykj8fNLgQdwn4YP1SQ/YX0
q1zN3oJaXF6mYzfzF6dkU4X8xDZBKxGjDmY+NZkHPElkOdnHma9HPgWuKVKGZXxV
ChYtpVBj2bn+M6ul8Q8ycPKtSMMELY8KmhiryF/yU99TU8XzDKnfMiRfkxXW1CLI
YOsCCNj88VMZNiqbXkbJK3ttqnyD0HtyVXr3k74V223EszoUfaU3bjp5M7mbQVRe
uqaUkt9tR9Vl2fDGZO+GvQ==
`protect END_PROTECTED
