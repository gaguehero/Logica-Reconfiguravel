`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsdWNc9nrzZKguXa7Iy7VDfBp7+QJqcwIcC9wSd1nudyVybk5SI3i5xVWRWHINib
KDeYIBL57T3R8D+x7qnhxRzdhBytzE9oChuLhYExlZ3v2BcaS21I5vNe15n+qkIs
4Phz/J2c8g9g3wUqODxRtbV4ueVP8DgaGzz9crubtdPKjs3O+kt/uPdT7Flhivyc
6liry11bZoHd3IPV2FxCvpdsRlvJcOv1XAez3Y/H6GDgXnkxW6yiOZxxuGMAwIXW
WJ6bn0RMOPmfdbBIDyER10Ox+w4D9ZF9oDvSABTCsyK6Aza9JQCIDTiCuo2PJPoE
jJe3p7t4Qt1p0DWUIMqXIVK87lc2amazuETQSIe4H6AGa36ISmB1RLOT0SiuOQob
itD8yr5cw49Im3RTkdqmtFcZBwgNAjo5cXLdbp8m+Txj76QpMOsGwwxY26yRNBBo
be5qd3IYuGwMVYMyuLZbUgfV16q07sRxI3mtmLVUHTz1QewJVJREhpG0GWQlp9Uw
yRgO0VpKHVjbu8NA2wOkM4tDTRD2u2SDAVHJEjY+2RDle3f8XOlWsIPlS9DpYhk1
gsnG0sFPZAxW4tl3Zt+4ZqrSqcbTNikWy0MYACU0e1Ij0wFN/Z+2oEaOGLZHn3e7
C5nyYA62N/r+M/CmqaoCzVRuP3NowMr/uHyZR9WE3HngS6KplBGSnDAN9bHQsX0v
X/zRD26kFajujBugmLFSEQumBPP4OGcDbcNnRY/r7qMcwvtAML1MibgVKNuBH65g
DWMS0Fpr6mEfiH1uoihtgwSSVd8ABMs7lGIjrFCjOHkLAi5IrHgaaJBOjRIYYghN
CBdPBUPz5h6MQBWwXOTsgPC+ECNQ6JyDtcC8umpqOpizVXEntwLrb70YFKJnze33
SnrvwrQkL6Okz4uPXZPQrXWzQjUperBvhDMjWb4OeVHdynN1/OVzJsbMqWxPxHD+
38qsapGJAO5BIIZTpBuxsSnU3yjHzRXlUX5gsZRTxJWZXXGdXgVSqtATKRruyzah
ZOBhqQkdhp/DipvwUwIxdEP5J+LjrOpe8QKcxPwub5EW+osJNlbHJZ0YFuvieJLr
JBIEbqc2wLCbLzNynfALSlFWFAUdM7/HujA3hMwZez2fF4PF/EwZODuCEAzPysR2
76FAhs3VLBtEi2cHu/lfyNLpcDb8VVBu+itZnH/5L9kfO1tdSGJNK4hnr4dEb/Pl
LTM+IsArg4rpvWupuIyaYrDvo1zVGjidNHHNhSkaZuEMBr+ZiODaaqdWOBy9qIAF
apqZc2g2KNjTEZ4jsx6DE8ngX56H7n3FlCNBSIRhHTnHg63AcsHCCt0qZ0s2iQFD
UO7ADGHRJ43ua07MAScTQ7AuL6RghmcFODjKKCYdoYBRl35ss9raDNqB1fyA+xbc
xW2T3v4XR9EOuC3aeB94bUr2xzatGY4+rP8FzMHpa8ZzAmnR0YmngvyDj8I1IUPs
+vC1DbAgdZ9qkq6PjClnhF5U+OKaXdTY7hn0vF1JrV2ie75StxcOkdd4FQXKVyOy
d7YDGTFPjr0VqAICGnnstdr9MgsPpG+Tj49QI8VHpKFutiXwSB1r+IDy2jyleCv7
6MB66Uzw6u+evuUGwmFVjQBhJhWvzOTarGl3cdC5WFsQLypQd7/a8uU0VghQphCX
xMW79/N6Z1ockEkzuanSjU3xbS4VEg9kuXfqOAuSRtkAiO9cVdYiE8GIv+0dTL1q
/RISoRYZ35LCFKDKVWWGyvk08IkC1VvrDYHYpfOn5njJx1ei96NIBVZj8GlDzjGE
+8Oj0kQpBi1imwIKoQCoGYUF8TrIV3Skde5UQh8Wpo/Xm5i4xlkGuo3xxGlYFSf0
tQfDEblaSka9pjfJzyzHFiAVA3/1WhxtLzfyFlwMTBqAB4Vn8NSFSTP9qEFf/0Bb
/jXIf8GQuK7yEh+PTzGE1rPdi9aXqphklgwzIUQWu6EiARtiUtyJOo3X6W68f5HA
o7mY7pgs5IpoIp2yEBlK8igihSnvA2iHYB0y7cO9HLA7I+EASgrLCMwbrGXtWTyh
`protect END_PROTECTED
