`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJ8wIGOes7xCvBSmCwGHt5Syub/KlPSg9WBKojq30EEluibtdcYbKzka/v0EA0ZD
qYyYoNSEaY7Nbh000HOKgD9EiiYkCJrqvkYB2HM1asxowwmg0kLxsEfSrteU25y9
VIUHTJqLuQs8D2rUq/D7edguWpixcXPldrb1iKiFThnsPg2Zfng138pYmBpTC3iG
LhcAPemPf0zEUUj9uMblzOw0AIp59YIiLAjQh1Xg95iv3Db0ac/Fc3rEFAtz3K49
UeISOs5XseqMDnPnLcThUjYH31oky4UsPPJuPotTrtPKcGB8JEAoX4Qt7702eY9N
Vwc4oDtF+a6agA79LOQxl5FapWooawmnqFoRWEsnbmwE5CDdfMFVLvMy54y34qAA
ekfsgeeXo//dhw1x08lScs+Il7/caTKJHkbUWGvsoFsvX005gvlidqwJmaYe5Aen
RCmEqB1zTgrDwpa/mDcGx0Jm8VdpNOsL/UPbctU0SlqigrIUAfr5wcE+LtHXtyN5
ZZuD46uno/6tFPB9uQYNth+dDx+wYxhWXLofJ44tV6ZBJIQcrLSVD4kCPDGJfrrQ
aqQaGxXJxGOcScH7i+/FRN07q4nzo/fDxIBah1RzEYaO8j4Hj++oy9AMIstf7W3P
aO9Mt+/+u+VMrkaeyNihIlK8ceYujVV1mLbyx+73kRMy2OtslIZEoljki5Td6iEn
`protect END_PROTECTED
