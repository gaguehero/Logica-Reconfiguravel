library verilog;
use verilog.vl_types.all;
entity totalV_vlg_vec_tst is
end totalV_vlg_vec_tst;
