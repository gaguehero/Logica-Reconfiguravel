`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7vsaqy8sOUjyTAomQMGaMh1Mi0MIymUhrgk5wxK+k8ntbDAUXiVBnQl5flkogVJ
obq6tQ8qnj20iSiYlxaHFVL73CAXpcrhs8SnVlDAdOCEVujUEvvEsvTBfvPXJNug
7+lG1s2siSxV3ybhTqYULf8HWzOrBpf0tyDx7puDX91CZXEqLg4MLqMUSr4n61dX
tckZhO2DDbm0vPNEqAHYfxQrbDK7FADSzueSBUCiLAqbKc6xXVjdCXMV8xqmXjr8
55f+HH/MeNvSg5yur0ziltg0VfwkMrXfoUhEtjrs3k/5PntGkoNItQAthgZsEiLJ
AImPpkJ0VwZuwKDCAHVr+3+zbrhO0xuQMwwDlpWBIDMCRBqmswfFJX4jHK2oFuMY
1klcwNjfk5bQilMMyvwEDO2Bqyhxjd0/kNhX3l0FWE+o/2kU/z7zwITY7Dz5dEM2
EcTETWkrtr/dvk5PyvH6r0qfZhxyI1bsbmkEGmF/3wQKMWL+LfuuZfV4vE0hDffh
ksRzTjHJmbN9MnrkRSo44hIlknPCq5tYmvzTlhQAbmhHU2xZgFR/qHQZ/I6mroQH
/ZecrrJ8okZtHM0Ckp4FvVNPkrGfXB9/zUMpXV5IJ6l2aUqVc4cQkE4casgdaFIf
wE6V+RSBBPXYIZhC5fDu0H1RxIrk4Sdrs9Hc6oDTRZaPSDIXyH1M/MUll9+oVmR/
KuHORXoaF2YhKI42+vH+Jr54V+Es3m3teNr4WsywzOaoKbHjZyk8smFCY5HDnb0x
8PrKQtoC+BPTONE53XsoTyZuPtv4v08jDFP7bO/li+sLdD/9E7yW7kZUeWcMDpdP
Istf50l7BXKV8hyj+VsyoFN6JMbm1uXVg1LI2u1aJG92BP4Z8SuYLggNxUfbk7fX
R3B97kAyyLm+RB0gqX4N9z0+jptMSKsJEi5wKg+SF6qa+Rg+g4/lGnebvpSley0O
5cZ/iV4GJ9PpetOd57KArkf+Yx8Tc2+QiRsInzscIUXhAhPXj9jeASu1auCoM8Lx
rebeagjVdzSzh3p4bIWBIZigcPuiobdq1Lu6229IQkSu1LCq+rPGpvV4COkIR9Hk
KsfcjVaizeIf6sonx81klbNPeaVVANDQkm08HV7lAu9nLENkSqRRrkR2Y2eZ89bv
N2MAXweV/iYBFYHwBsQ91MDzWjjRBvRWGEb95uVlv6qEiYMg7bja2Bqvaf9deMnf
8KrTAy/JuYXreNE9bWG6t9GkDGRo+QE+VAwVwU8RVH1EMtbbMzCeOSYTV2N0tl4n
OURQustFMDLuXQWEFmWgz1eL6tpxaK58o+5bHO7sXkA0yrmmdkvbbUH6Ye3TOz3q
7YBpAvs5NeeCEZKY93OYePzdKXbF03/BBIPn9Q5CpZTd1/ID3SwqkhVuL8NaZP8v
Xt2EzAP87C0TXifO7R3tGQuR+fjKx20XrroxPghlcUPfSETrRVCCbafmrkg1ClaF
RQCJPHbtJDYH1WccV/h94xXXDQfyy6tKQ/bP8YPg3/Z6I3GX7n7bRjqh1Shef3j7
WvvDNRBDOtumNBobeVS+PG+YAe9jp08t0y6iWqhweEZKGCByEonPNph8HWTwEosz
4QUp7vQTOFuR3zfZfV/CyUaQuAP05DIXsloqh1qYSWqihhS0xNLhtAWu0fJvlc5I
zFtAsvNoWtN7V+OavjTg7w4tKJ6xwX/vZ4UJFjutcyDwUD+DTm33Qvm8pw3STbE/
ymgBVt6hTJcdjISwoZTCTmHu9xN2BfO35Jie7pG85UDHncl1wQ8ObeMcWvgcgeTN
L1y8el8TK98qY/dUYMVQLL/mW36UWEJl4LDdtjKQSgPQws/2zi+XUlZshzE/wydS
w0jwk0RrVTfTlHqlvqHBKLQNOLv5Ixv9ODOQRU9MzBzCeiMGb0ltACZmY2dWfqUg
wUmoMTLNhMoqzrIjQAU2a9MEIy2EKwzsvh9BxOFVkdUOFiKZ2N9otocf4Hf2TvOR
16GytfhxsfdDpwHI6+es57V9SzfdyB1PJodUrYnIXMm7CZykZ7YpOBcTxLdFZgv/
gU25yl0JJ1PNFxSk9+gFaApnb+vRoNucZg++/4tqmBAtLPVSxPFA4iEuBDPippAI
AKdMk0VNk+iJHalEKwH5kb39/6Sxf5uAMwf9f57CXDKPtFBU53XYSZzTNfim4svn
6EGxGnykYy/h85hrLeABYmqwG+aVhzG0cO3bkzjNrCFH1K7ZmkIrD0gk0v16rI0s
+0e8YH6N1nbfi3nlVNI3xBPfuYkB5x7xEqr8pbG/5ZfBB62XoTSmXiJIplLfCw9g
mRZAlkjo4mT7KTAkTJCoTLDlNyYlXL6Df15lIO1k9a4DE0Q+c4UUaNlFTFb4cOQy
ZceE6F71uTVHf5RS1grRiJ2rl8qTdHPrfGbhO9znJ8ohA46631s+v4faEdLlUAOt
QSX9v65OzU4ne/KZxSJ7eYaS1A3bJAqIOdvD9yN3Fq30Hrd8StBkl7Yje1D4Y3Vi
ROgzeGaD3ZX4Xx0NJywQKGG+dvTUTWUbwQbqp8+fgxskeXob26U6xN5Eysb+4VG8
dMBiNMOXdvAi6ecE6ga7EN46AScXW43oCW4UJXpJ86ki904u0aFWq5x/VXz9UECh
KMH+tjxvSVjCe6B2wF7UT6DbPDevSfRVIUIVQxfcjb4q4e7O7osDdKXZrIO7gum/
ngltRhRc6H8nfZAD3SnyBPSQKYqAj+51NxTJzTqXRrf36RlHI0jODBEx2ann4LIL
baAA6kkPhnddqDLAX4RtSnnJMhP1oy5FHqhnhg4533JJAsKlemQZH+IxeTry23PJ
J4pSa7ToeF4bbjc94dcnUxYMuM99bE5eUHNU8y1kJDxBRc2brP1nxVjzzHRhkb2z
7GRBr2txmQU9Y2h4ecj8bM0PLiBwWobtMDfdARJQu5Y3d0wmpLDoEBecHr9ofsqT
RmqmdaMFiHG1ZPajFBYoUdb6XpevJ9piPiLBsH7XdMkaukLLAL2kmGUjbAN0uiQh
QE37G+SlhI/NJPjPFldXUyY/iMga4gtEiLjk5tqetIdgsVImH8jQ0NNRugyG3ooa
wh8cU0aZtO4bpeWcui/eGoIO54zUL6Cq7S1YvSyfgBPHxguYd9ONjZEDEx33aJos
HfoJTs8RI0mbVYrWz9r2rkfLPfJGipqDyOhlawLDqeQEwBi1+MlzbSKLEjh3hixK
dyZMyVxa0Ixn12IHEqRPdbeaMuKF0E7ct4gs13+0q48oPQ6iW8nIbmCU/mKuoDS2
XcQ03DkYwN7a/zs1KebAJ7GnCiQPvMPOMR37ZLHOA9qNTB4cLdWrwhUaqpPqSnR5
0Pazqs/uAsOGw0xVh+vCCrsmf7RksW8Q//lT3abfEtcn98zA0aSfgQmQBMxsKWHp
WDXTjgIK6njpa/hiKr5NYaOjs+DkF64Em1VOiBixOgKVY2RvrPzdtYJ8yIyP7zQ4
yVp/pySxMEYlUCbreUGmQUify0CEt6a6ci7Z/RKyz0ZWPnyb0iQCjuObZU/KzqRh
V2JM8oKc9NbFpsDp4u3AP2Vj3u8Vt5MdsZQG09/4/zVeZBTBM5Q3agft/64N5Yya
h6mxps5+TL/w0h7D6Pz4LudOVxrA7X8Xw8nwtwZkAYUaC9nmpifY4RKhk15Yiiqf
gQnyU1tP1pKDzbHOITQaNWftF0G6OddqgZ1urgPW3waugHyElEBML9Gkd4xOzdNj
5e129JmMh0Z7bkAONfjQq2ID2kDo3FiJtHxLwBWRPc26riyaR5k3j0vHVIjG33Gh
lXsKIP5CFeQEzhgeffGS11Rd9RntXTfLyYdyfb8UYXxmD053Az+Lhuuzdts08Y1g
HMyYv/WtFWmMVtiTHmu2DGBLSNlBjc2oYZlEiAkYhcLeZRKYOUVtNnf2Et9zg8Xw
arS/VIQEc67JBa0YCAa6fCGq4Qmd9HDS28evXwTOYrqkUSSZp5tBGtWYnaRoW7Mq
1DjPBDjIpaBEEk+5Ok5B41oVOZGVrIxFKuHrPQrrSbqiX80kXPbm2t7fF3P9qFvy
oOlZRuS53kSi9T8c+gwdH3ZmRq06rUUl5AWI6dubustBUCxF917NRE8cLhKJkhEN
Vb7kOGeceWdUjC1Be4CZ9NtrozYIu3I3qalLiEmlLziULEUCujuaJgmacXOz6PvC
lRMNCz3ZMwBm2unrD6NWITiP/VEAbAd5lTgUD/f/KbEGG7sJVw5yDVaN0UYI2PAn
FL5LLRThFYW6xXxUW1rk1+0PJxmt9nqbQ/8w0zSy1sCD6R26z9Mx3MRi+75H07iA
Bdd7Zi/U7iMs/30Ehi9x6EaLptZl2IEVQCeE+yi4rZXK4GgsHdfEY1No1hTV5ch0
NDsRFGbrO4m6UND8enubl3KtpUCzUh0EzLM+54CjgCeb087d8pzCP1ErZuU+bnfa
/Il0jvaNH32Kwowxa41wKXDl9z7H6qdA4PZG1U1CqB64vQPu9GD4gCIYpFhaENq6
Ly12KRwKqOYBCfKapVHc8jJiVEOkdvrqHJWxN9MV+8nZZIG9P3H90RTiQMkvTKsD
GOBvL4nNAefiazse2vCQoVKQS9nvib6lcRw/nxaEXyNWOPmRk6Na3UkQ4RjD7e64
gASyV52vSWTe/OF0Bch5UTG2C2OgzSQY5QZe4rgJf6HdmkFSuBPRsBow/VfvJBD6
R93K/Kb10fJwBQHhNXp7WhZXkV80+Nn/z/frDy+/6vlgrPPpg8MUjz+XNdbGgytd
4KYBc8BJMOZLSjs2b5tqnWG5jlYsKjkyh2yuk26MbkixGf3ijngLCESEwlEYmZ5J
/caYlz4TjhcYMiWoPVewrTYcXenU7BtBKmYZLrlKVZGm7uiOhJNW8ON9NFpi3tKp
qqMSnUEKkV3F3G/Ui0VQCA4saqtOmvMWKAQf56GF7EzOSTyIQXbtvRSSk0tdnSRC
6GGxAkwjfeQzgCcZ4T5PczwiuJIZ5h4GC0AMFPYsZF+scADmPDLDsKbhopi/0pf2
oedYfsOw4P6x0wQEx3/fAG3Pmjs/fGPT2WKGNTOMvJYDeOjjDipkSKkqvVuAMCWG
DgNOJLSmm+1XXqNZ8Acc4C7gCkS9Aa7/vxMsVVxpEBfsLA05IauR6A6gpST/flbe
KLWM769MHlXaY7hC+MOG1BlVusvaAIDJDdY7WQUfCnhAXk7g3psZrZw9tgh62lVg
KwLp9/AniNreps/SKfe9kg1+Llse5AfsU1jgejg2+lTG40XYJSZvM+pwBqdbf8N+
Dl7HB2CkVkLg6aw000xhe+YJHR6N7gGEcZV4vFf4KWkucj5Ur/zOh2KUhGHR8xFG
R6aRvWEvAN516ZIdmf0t/Vns1496bGq4dngpVq0MYtVzhysBC+PpXwV4mT5CGBD3
kpg2phMWly6Nb6Fekyj1nEKKKWpxDoRfe7Rl00jMjTrhtxD7DGWeB1gq3z0dVZTc
/JSi+pvl5MsAkEXdUV9HWLycF4aFwblCRhBDJA8AqFwtL2uw7mjtBcXu+essyqnN
6TmskyuriwJN74J4H0PAjA==
`protect END_PROTECTED
