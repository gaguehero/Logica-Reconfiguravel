`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XKwdqOhqJamK/255t8umUGqXqx2FdBOh+GIq+4MtgojWR/ejTNQGcWKU5y6aYB3
XcZvXnO8VasAN2vQGKKg5KrTuaqaFOJZw8cSgJ8YLAMNCPDXkdF0n57OmONFNtyY
AA240sr5N3emALEsq5TuKOPDEauSh81Z+GC5ZRAKbhh6ZDX0a7ONGe3JWZAynl4S
TMzEmgRnejhCQtu7hNPXxqJdeMJJPkpAReCSpIah4a1Zmoc7Bnl3fl902xbSHPES
/Ch9YTGIVHFL+tPMWcPriHsA8pmGO1DoJckz2h9pZO+qWDwijEDUqZbd15DF+X2x
1dGMVmb5WBg5eKvrnD/Z4FwF4GV7wcWTqbG8o9pfuh/OAlp3kxxs2Dk/YdkfcANQ
jQFDWYLFPmS2y9YX/EMe2KM2QxPl2ZEW9hagsKT/p/y62wEj/BPRNIgvJoNIqo6s
Kp5QSc3INncPoYBMT/KfUJ8joELeQi/z4wg0bl4Z9o1K2nq3qKJtGyER/0EUjfo7
JTD7JWkB3nVXlhbaJ4/hj/EaIBXS6P5H1oumim1KFJjRsOcnZY9pP+uwyZmFxVKo
Ikiv8+UBhMNSdii0mBmUpXqQS5DesnKOVRo+fVRAYdVtdpb7kBVvU0SvlCUVKpir
roIWjBxQbR/6GscujmvyCfavxtA6lkUaqfIweu/BPsTvioez73aSZeXWfCVMht4c
JwUVAfQ+4Wzygy24JfOwSPc8KIkRa6/jOPMe0yhomZseK5YSJ8w+lpInrNaNlfmV
hTXAcWlgyjwnGQagAL51+0zPoTCDUdcteYvIbkqppBrGZcfmsxlovnKyWerpdSGL
fmemU5SO3QaDQR2as5CKGrq1sojRUfEzJlU++D+5utnc6CK0Ht1+rfnN23R+DFvj
JKeNfmM03uJGhL6TZ/x2d+ov+PNjWMRMts5IzOidbc172tk5Nu9k3fdIkD02/1kU
rb2p41jLFpsVRwnzH/mrSG9h1TpiMDhSHyQFMTVAhOSqhIBO86UsX5AOh/j4k+ki
ErYJZjyqTHG72o1XoV+vfe2/uWG57erhHjap5Cz3wHEGm92YwE58bW+SqFav3evT
IT1dk/p0pRsxg5Ts+O0n7ZkoZn1Ntj+22AZdLvd7Ort7iGZPUkZycSzOY93b9npm
g35naw/i+Uz1H0XOLJ6yXLj5Td1lRhrmbBrOX7HDuzLXbst9thRscnXwH5xyFBq3
oHMD+5t9C9Ud3Wgjs0pBF22VAqlU+gyXiFA/6BUTUKs=
`protect END_PROTECTED
