`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oq3r6EgfDbBE8xE5Cm8uaNE4zK1udRugKMXmjtXdNS7bcnYO9SoQ1w/PikdooDla
QuZRRwmuy6xo5WxvHYCBmSBXn+Tp/Hf2T83uz3As+jabnu9G5aP01yel/NSZWe+Y
7bv+yN5361dTqi3ieuyAT4ijJKKcXx8wiTM8qMtHgvxK3TGhCnvBSu7PEluRAwq6
GAmMKtDqAUgeHYymTUG1ZcTmI67NAmuS81FUQCg9F4XCirO80HqERO6x7vUHOCh0
yeepuKK3eXX6IMsltBn336NZzo1iYcXwNuBxlldou1os9+x7qxRFUsdVVEELUFPF
EVjsFkUK3hLPB6MyOSSxJlUS7m1icU8+5SJwafofS+vTwwLkaiMzp+vMVNjEyKcs
jifL5GgHxl24hJuVr55ZBlIKedw41fWElsG4y3Sc+h8HdmYK09obBKlvwu33gqUI
Et2uH/3mpFH23Ib/S4TYoSnZiMniYY9OnkDvZUeM3rAWWXgpVsDEzmma12jiJPxO
pt3G9q94xP0zrtT6X+A04u7ff13SMWvS18vXmdS10J/s9GsrMGvfd0bCzeIGJqj1
rI0M0bLf0KgVsbJv+VzNHx2h+oEYLYzJrWFulqB0dVbqt4gHDPXW7Qd148MN0jIN
kTq6ltpB/+THltD6CmVIbw==
`protect END_PROTECTED
