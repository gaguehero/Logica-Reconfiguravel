`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPR2EXVH3SJvmZIPcyjK4bg++NBQbjjJzdJRMfwzfZhkkw9hs2XmM4Mh7nveA1H/
9SbIIcfs1nto3Ncaob1Dc44f0Aw/OpGLPwPvd9yZpJtj11ZuNmugYrOGv1ksFmlr
2V7iRTVliXDq5vScHHdB2lDeOylnTx7yg1Lxzs1LzKM0cbrqBp2YRkrmB8qnA5N2
09VN+PcOsRpw/YAr72k216LGgUs1WIY2arlzbHiqXfbNOiuZlNkPa2txIlpXy5CM
bLMp9LNoroLONgIjl3bJyMxMGnrCrwADybDjq2ZmVLjOOA4F2yGwhCqUalr+dJHq
RZYbV+xCPoyfiobzPLRAJF30dSCBCZcIvt0ROit4SPuNG0GFNkBfTsz23Ju8Uvy7
Krr0DHycjwDdG6+BlBxpP1osByuh/z35rqCwOygPartBQsj+Mbumtz+uLBwn9Zws
LVb/pSEliWkgupkG6cj2+lWSPqxOlnL55RlEATmI5eQi+8BT5HSuHaS/9/2Rnyh9
YrJ2j15SiDly3+uiqbNHMpsD7q9xCQs3evnwNYyiw3oYd5SETDElXBziVGBnpl3m
0mckTkvWsCTJYfvB+VU6eI4/3FUJf4xwa66if+bQxQTKtbu9J/buqBF7Z3Ik0+li
t/C1uVq5nzvz8iCBY9VHh5ZurjeipZ1JwBDGV5i4rDbhRoJWp1FEPJ/+R4LcEs2Y
eMDFauxWse9uGeZ7ocbALkgL7oZoblaInorcXSzALT9Cynvmytez5d/61eoUvcsy
Ws933pgvu8Q/NmmfdXAElsIU8dMy9DVWPmBVzHd8i4AuxwCrpYx9DrLZWmraU3Rf
Ng8FjwI0y4rPI8MAiTQiJ3NuqMkwPYKtqTKJF3secCC0qYWI9cYkYAQOME+wdghA
Ok52RWMUH5wNftAGFgz0BV6TFRYRJ65tVsZ64ogJ54I1egs5hatLq+NLL6K4C3Dr
k70aeZvZzEX8c99YfsrDbeS9Dc7/laHLgJktwR15VKyMRJd4pLytPohfHBOJy+eL
CoLZuojpqJWl/s4SAQeiUcxYXYnp1o2pyNH+H8e4cOlKoCfKNGjKJLF2TDRQqHB+
qL8YusClRl9di6q84ReWzvFdiClEgdmsDIu0D+lKjArz83VqgzltarDlPJHjVV4s
l+yINyQfGoGiHSbLufk2J/m3vd/m7D7o2TJt3jTRQHCn2F/rKtiNDHGUFBIspRhh
lle5KRsbYumKyQJQuEjg1vqmTJhJ5EJouTHM3RSA4d+kinLTej9JGbQMhSgXKnOW
fNc4BcQmMjS8BxuJ9qwRd1Swf8O73j4dooH9ICBumMi/WEwDyzKMaiMzx9bokjqO
2JTIIdOLVniZQfWJmSZrMoyol76HHQAxyQL7swD62rV4baTKdQlrIAiNlRPf6sNS
FJMWfqvXSk91Upbm7Bq6AM8x+UC69Ty1G3CBrOvf9hwmr/23wXvGOtkJYhoVxJjw
8C7JQrVX3tPjeyVGF1enu0FwSH64mI14G1l4Twhf5JCv0MqG4AdHi4UEYNjV1lf5
SdJnbaDY5+zdiphM6C2nly2sz/SjyATfrYEPOkb/xeBIMjm6E1FX4+rEFOfLG4Ap
zE7mD8EzBiVZJP53p2riolUyPEYZMrleAAaxg8brepMcyTNPgeKSWsgT/r1/1xR/
pUJRPAAz5e1qWJ7TYkQolvBgss29egEmLYYOz40lSSfl9Pft8sYbEuvcpa5orEwk
yVnkEB5R5txJUYRRDe31AbIdmO3AzXotE84RuBRJLIZipH7Rd7eifqHUZBMXuc1A
EDzARyGBXDqGbYEYGARHC8D8QnvosY0rXDZTY5KKqh6HnkvIWAfroz5xdSPd9exz
72IKQ+iRB5IKWIIlkC4SD73rJxuRXTlfITSkSq3T9qylD0B8BtwhLKajHpMaYFe4
rexiJEf2j13nyC9XYNBZy3QDzZJiDG3W97C2DolEQLvvTsW8EggwRFY9cNrfQDP2
CSdsAkHhLV6RUvQCOxTSapPNKkFGB7rCILpJT52MlgdJz+uEKeJgy7X0BNVT0fa6
fqZboxFwO06QLfB/E+4flS+jC+UYoKC7Uc7cXZU7wK3d8fofGSuJO0OnIxgNo+/p
65j2M5IejRyTFCiQoOYfDLfvsYjHAIuHFgUUe7b70PwM278B+hVQrjR8hgQEW1SA
o+4cTdqs4yS+vz2GWp79xsdIaY7tbgfaHD6nJXmyAgRO/pByABy3HkwbZSIQv8q7
Z9H/OJ4hU8SrLtBwK2YfRWTRTUj3E78bIFQRPk6ZNG8A4FehW3n7CXvpcDiKCdjW
6xt/52aDy+gE8bnqG4VZqClq/Ss+r6nvhdmUFOHVzPTvUlynrFhTAkXv5TuA1vN8
t5EmdYyChHUBkrtU1xCiYpyy3h8ELpyV8QhB7I53RigOacZGzOtQsjEbK7s8NvSt
9h1JQocsfOVVjckHQaf+BYpMQlOv3RkI+Ra5Hjom2Yidv8MfFOjudLMtnDW0EtXY
IOrgsvp15HjR9hBqCHb/+FR8CzVQqFEcFbXJd1Kj1M/WmJE1qr/vxKUqOfCh4Y2A
vBc8H3K53mNXvx77FPIgCPeBVHFeLJJYAptHIdBYCzUNZ/bMD8xFFhGazWkVW4CS
KSMnXQCXAZprGTHaaAA3N44FMcbaSL3cwKJ5JseovQAwyOU5L0EMmY4jnzGWCYfH
r8oVxupu/rmcP8IN27w08yJnCQF9YRTsdZFfrjCVRzneSvLYQMUK13mRA4KviV9b
/Q2FgQMMnqGMcEgYA4amtSD0FY137JRKr623tYRWTLbXLVNsbEApL5TjvWqxaVft
cRXwhwT/XUFj5ctvwtn77m91paqZIS1kaz+IZGCUAM0VwmdY5X5mCS5VbpAHYNPz
MnA/W6AqGKIrHy9MHQRijOD7y40ijEBmTIu9MnZfIJMiofhp0mR+dTipwwe0DI/V
AmFjjkl0cYehiUiIkSN9KBty4s+C0FEpioiUkpNOWGrn/KqCr9+Y4J0sBQfvLwzN
81YjqUC/OqUFHgG4G+tqYygLUS/6s8vtu4VSyhGMbeEEI27SYcy8kzb0PJDd9+r2
pDim0qZQpXv8DBMMwqo4o19m5QsVaE3FqAYcuI0zJZdKVpI27/ugXCGj6eygTbxN
7NSYTU9r2OZ1GlNNxwVgPlndVsAqU0wFAf8i0Y9IplTXY+1XzSss5orzKlSuw3wg
Mn8NoniylxG2yzkDiJ3QIenanrpJq/quqWEu1BFeW0LNisV2pkmjJ+S09W6LTuWs
8ifniDIBg3MvWOwNTEeV+3RYm6JCcII5RZIsbov5X519zn96sLsD5FhrRSCb6pyW
yQz14/nPmxI99b2IAQ+uhgsx8WCH9aZrlwD9lppXo2iykIPGTT/z8uSMuEDaVjBP
V47q9LQQYnogyPttJh62V3TEUXukBp7Ek4AYdN42wmWbhU+rL336O/LubENiovC0
n8H/EKaVMfJktjrpt8cZ58aQFLibsbsAYEL7+whjmP1+FTfzf01vXojH3SrOGwub
uB4+k1FQ22PBoLz7Dm+UphJc5KrJeZWQatdRfh3Wg7kyffl5WMoJCXxRmdYCSYG7
u89OGuDlW9Ge2TTQ76bghIExhMUkOVOhN3/KytUlgrHY79tDlPuuXn32uCUANnIz
3sXZ+r9szICeEfj2IFnHwajsehFzRAfrMx6/UUFBgwVdkWcbXgWw/Qc0ezciegSL
7QEsjWb7DDFpUPSaT8IAzA/oYwx2hdPRLRXlQDvuPewdp6uI7Rwm3GCAypoogKHf
MjvR4dYamV/f1tTUcNTqkMrukR3xwxbVYjtLhKVDEzWEe9Ds31jJRIecWjHWQaq/
RUrUDWZETiOO6Mi+83MrSpmgJDP6e+wS0d0Jt/nABLx7whL9bPNrTWebbVk9kmSV
/PXRcWnhQrg9DeWUouXueUcTiXl/r4ApIpyWVCJSCUhf4OoJAJWLfgFXsVkYYyIO
aLFGHqH0OjXOhYxzA2bljVcLJDTFiTiAVPaP74lYy+U9KfRDjnf1u2dhTe2VEuEa
TXM1Jn86/9vcKiszTmRlKmwmErjVg7PZPEuKqCpEDcbsBtljZ9DKbpYLbDIGIX4R
ApKGFSDPFDUeeoteYNX53tRHB5rB86UO8crB9Na6ljH9gktM/LS7Yc4xMEnMoFCG
dMZxqRpkySUc71DtgXb7RQp+xjhJmDosPqNcO2GK8TdssKm3dpS8cRjgOQ7NbxAm
4v8qffVrvfjHfVx0bjxSeicvjlXb0ZFWcdTTsrlRM8L79vZ/8Hv28CVDl5tNXUMs
XQHcrIgrSBrdWkj0cvvVuWCrk829WvgvvZRguQJLP/ifw/NMHyGRvd4O5IEILKhO
4G3urf8wO5kBNs92uwag0GZqD16bGkQRV6d5/6McYgV6BXc7CcZccWD2DoL/LRUP
KnCONzPHeFgoLstutT0UWyQoGFr15NgMXRtBtC5BxIDOaYDGgvO4GGkg5olEiVYC
SRrLXAs8Eynp9CVI2fyj8AkZTpNvXXgZD5vdyDuWwxc8gYBwhmhh6huDfKH4XOnd
rUSpnbqy2rMBE4AIpO9RGFNkasJLyrZ663a92tVendZj38d40A6rMdKtdruJ8fkq
+yr8jadXQCGccJJBghcnpAxwe3nD9dsy2ZPvw0tXyKvwalkh/19eDiDgzO+dfB/W
4Qg9P8VDdEg3eD6Cub6pnT/QHcmkoITA2e5xsp0R1GneehpztCkOKWXSdteadUUX
uRAZaRCwzb7YHjQa1EuLgph7z9Jr4Bf7RIBEUWsdIu2aj+ZlpJHZFR7SbRq/zeXZ
do4YGya3NRAj3JsR264wwYC5jMqQ5iZCzF/jzbq/mDll5uH7g+teB6I6QW/m1keF
iQRIHsh1p8mC+Hk9WdjbRUIwVULkfBgzP56cH3YihtBohukMygrugwXqfV1VNHoB
xzAlPrJ6z1S+YiEJHBRcaTjPvr3QEOSEIxeNj5PLCVy2jrenH6xYD15XaJ5Lj2Zk
5OJgZ9VywbwPOhLj9KgvMVNnOw1pRUMFr4GVROSW7f5yldZIv5wZtzEKUjjnQGYg
R9nSo5oxU8sf2Ljk/6IdnxZP/HqWY1LcboSpY1oktKoV/q1TV2fcVuLg1UnzHSU3
oYA0VmWdYwPvYJ7z4L79j5lD0pDcgBNYsLNVkqLPOHv5jbLECIMTutvYqJsokP38
GTyNda7o6AvPtxuvSZQJsCymIUQNlpzXnl6K0tZdu0EaXaCUIrr9XKSsJ3SBH6Ql
lwj9zwoqDPuub+fnp/UOvHCMlgtjA29kXz8uNSu4SEETfkrWYaGhQinXMZ2JPCFX
/hyP05yunB21agC8MAvpzD1+7iNWNWJnd4UVzcZFDNYpnM55WLfGr42Kmyox1z/a
xKtA9fgqOt4qVCC1SnGw3vrnCft9afodVr+GUJ1n4fh40q4fu2fwq/Us5t0vmeoV
vi7tEQp3s0qz0n8yL4hUGtEpIJZZJJ3Q/I4crBbGPTgHJYjFCTkw7RJt1fNGKM+P
qwNQ3SGds6JTE9O89YhlBjw2bPpLEJBro4ZESkFpdrdPmVFUcklguD0Wyv7Av+LA
ZEslEOXOjaVQKPfhpHNitnd4pFXUf4C4e95PSdpyLJLkPOfc0Pjf4kREnHg59FSf
4e+bz0d0MmMYxlIJih0Hb7DR430lWWbI1/NnsBsOWcqv6F8Oy7Sfu4T56lW/1twN
fcqyhgAWAmpEWbV4tCVtfeeHC4qYCAJtZ5TTXqa4EMqNSSLi7yl9mDKvxPzd6I/r
4seUsujRtjqf33ZOUVMup4059pOiaHz+Z3uKLPNqbg7MbzRVvvAefw3UgRD7N34J
lGTlgkXTj9ZZ3HMfpJjY4aeNviRgyHCo+jXSqH7w0+NNOZqrjldPJ0SN9eyF+v51
BnGP7HT9VDgOQcBpkca6alweOd4z/L/85Hk8RDrv0O2z2dQf32Wyeh4Qbgn44284
TgRoXZgvYprBq292n6Xc4RhZZPZwjlnTAfKui4Wdvyb2lUwRu6II/TFpDlqoQt6H
HrnMrYP1YRbxIrH1GlBWIuJozuPPLlAbOvzimYucgCdzE2rPnKlgAzhKRzLIaO6C
GGnVpOsUDVqzUPQKKOOMuVsCDx96eEd3oyNEVv1s3OgADYvIBujuWJZbL1Otgh7e
Npq8jVknMmrYQe/IHtMCVMguTfJRqkMvSygQLmVOIof8dZ+NO2cuSBU5IewdHH8s
I3GiBrBbZgW3aI9nhJfDg7dffuE0jU2+SLMtemiA9FJKuKPnzlyV19a04rnQAqOP
HQYS8hMal7RpvZVm8AgS195t/dN9rjpmce+hlNeL1XVrGmuMBlRwaPlYQfRqpB4i
0b1jYHf2hoHHB8yp/lT70h4zE9uK2Gpu7iVtigAroax+SQWnpY51KY92qZhc2Fbq
iTcwXS8txOQD7dBduYwodrw/ioOyXvUGCURtE5yDc2Sv7qYooIhbeeWPUFSspb0t
m9ZnsRGX73FdtjpW+Nw34195yUq8iGcITfhkFSvZidYkqTE00ypxMSdMO/lRLdRm
oV1NVgwKWEaMKZ1O5fTbEfqgS76vYcNpy+GzNM0OvQWwDbczBWBoV9PGUrsqmv/W
DYCB6uTjRA7TMPmhJy7xYgnZzRmvsu+XG49JFmi32wjUhbOdfaLyjprzy7SR8mB0
Xay1Rr8qeAjvUUTvhvXTZFmGKbV/EfkBXs2hFkZNfKsyqfS5AnH4Y8Ocy4IEoqKd
IudTDog/4aid4F+XuxUHjbAIk7V24F3O5tVOGE3T7z4ODKi4vvuf1HORCfT+cgdp
Y2sRbdtaHeK76qN2LdMvroWYOMjF05yN7LsLfGVo7p70hixf/Xwkl3oeUj2Z5IQX
TCGH7TTdwZxLImRpnx9uuUNZ5kpFD1vVF1j7bit4B8z5RCy/ctYkl21EFHhiYich
Dc3Ll0Mch0nGgsvq8jdMz7Pw7zIOIe4aiVroqyZlM1dAHm+t4Xyg9zc+B7i0Vgm9
5pyK6EkC5ulthnz8qEkNsl5o4UWATCyg0y4mLzUmJOU5gK+h3hnLY5b2Xcj4WjRY
QZ5TfnA1p6NGX1L8SEbZqB5IZb27DO+zNxpan2uIB+w8kY5OfuCpH5RA/pOkgKWz
EpWgFW8IFc+Bssg/UkrhFKbJ/8eKW791GBTfpMZbXNdEl+T4FmI5rILlowAPRh5k
MWPmEXmdHUvhlUA1SautibLtMl/mi977S86vad6xI3yv66aG7y362MKHIrVMLr9U
pKNi5MLk+RXjuo5NpA1CsM9Gg0I/tvBvMVjYbBFh03qAJjX2plVi2BEyYZUPLYaE
lIiXBh5me7jY9YWVpVVGW+2a26XW7t0qwelvnSUyKozYW90CAom6Ef+GLD4VuIVT
+X/bSt4+AvVBp9EKl8MUkbxfYTrOUOcyu2VSQ8hfs8h14qgQixm1vNFJvWBOpZYe
0wVsoUqC2y1ker/6Iv+9wOqWJp+MgE2eyZER0Sx5SkzjNPr60DiS7EdJYGx7/O55
4McjrTA4HDaHM2eYRW88Y8p8mgKUK7Oz+jn0Gs4pFtzxT1BKulz/obrpmSo4eiIF
d67lBIFOnEYmfE7mM4Nnz7UWbEfazdPOrJWsrLYVYRukRJ4rPKNYW0Pj2K56Esa0
AjaSU0BmP8Lkv3yJ507+oHC+LQSU3oyd36SFrhfU4JHv21rPUOvDmC17CgQpU3gU
zFrhhMMy1Tb/8zkrFZ+FBJ4dUA/F1ehQKgE0TJN1MDXDEYYYMGfiabB4IsKaNtks
vR//t8x+8XgDoOX3RtIqehrtm60et/lY9+DQG+ZKVPHj6PIe8tQDAaFx5nqxEUw/
mppWw301QjnEX395klxAqAHMyQWBTPACHtVHnZTda3/y5ZCSf5V6bv4kxH9UQaeF
PLiGKmRW048AEs1Ep0Zs+p05EauYUpmpaq7oUlgjOnqNFxCTmdDzQkHZxO4SMrL+
d5U2KofSM/rFCO176G9BFjPMC3hy2qDy96jbZ+3yBewMB1/hvkl77RJrvkopvWmW
k5JZeMD2aNAPeR6FMKWcKSBzUTbviEOfrVTkKp3Nh77ANf8YM79DwjL7r+0ENGbH
MUwtqyP+/96LGZ6FAV/1dsaSu2J/QQptSUB58h1BJcOmtuwRRluM4T8KaHcb1xRp
IFjzpdVv4+Ie9+OcQdQJr1i2Rh4vbR9BqtIgmypchcDgSjnNE8ElfGGmiIik8nbT
Gajb9h+QvXK3dN4p1aFz41fQ+jc2aUeO1BWv/pGTTMIVGfaGUFxAIOmnFhRWgCIw
FPqVdr/LmccXwaWoPqEvoHZNIPeG3wzFAWxjJBr+ZAMPHxzYL+CAJOKR1M4Ijd4S
5QHb7T2dEqKLVagv8YYuV7QNEDle3cC/L8/My0HjdhyzXK3eFa4W6KfA0VKM5Ivm
Hz9QDyEh0bn2jJByY4VeXOVAFeAZ81cfrySj8KbtghvttlWIw9xfzvquSUoetLJK
4dy7JZHnSWTdIWh1WGvlnLlboEpuqbwcyLQm11A3Q5CpFrUm+316KVaLfIMKOqU5
Rvjw3rNSfT0Bvr8N+BuGdUVHzEhk/9AkhMxdg+UgXdgKH6i/pgSWW6Cqi1sLxkBb
46VRtHN5NKcNEbd8XbMiDC5JH2By+cU4JbeXTCaGrL85HHhbdC1cM7BHl4sM71+p
w1kuI0IrjAqj456bJYc28mi3YDmlm6fTnNn2FVWzAO7wfx27m3m7bmuxvK3qXh2h
sWBGIV1Va5dhRtuUKMtWbo1wHGg6mj23FdR60SYpml7FFdXQcDPF7gK4dlJtXtPq
nE8uI820HjgLXdYxtHTFpnfakjKawVQr3PaaQHVOR+h8B/9aV8I2rho+EQ1l/DGb
DlrHX/4e+r2mJ4oCuCqBvCd8i3UIdFMMzQc7tKRx3qU4QbkGMYGHrvBpdps3qtRS
wT6s6dsDoI37tuBxC70JnOVbPYdy14pUbdhIUGKVg5L6Qa8pS9/1Pn9atF9g2mZD
QDoFY8WNEPx0mIwhyQgaBjm3ArgZ3An6OLHn7+JJvPztY8BLOtSnMhjyuky/TrVo
9QOXjJ5XDkD5n0KgSRzzFIFTU+1OsWUAOODggQHX9WDjfaemGlNghKyNax6h8Ilg
uWrm3ZCtzzAVC5oltc3sYRIKBRxQVDj9xMu+Cw5GOzGVqt49ZSeOMe1ItWFPCXIy
MzylpGbS4gEiCiq9cescflKLnqkdCH9MsXk6Grg4SyBxEHbrDnxwPnAowWcEND+d
QyM2/+m6wWOSqeeIIr8wKO62BOQdA2/Yma5LzI9HKjILvcwnzaz+nLCd7J0Y/7h3
NQHolt1WiEOVVtTG+7CLQ6QjK7m1z4fQoL83BlZNrGrIXpk7hsQSamat/zknIW9l
+lHcy3M+RRmmqScYYt42+LpW2caXA41dIq4ReuC1KkM7IFVPH17NNRaB1tQzaZXD
LlQNaYziAo4FS1CilQ5grv3GHIMVy0gxHMx2t5eFRoknuUKesYUC6jhR26dQ+E5d
9NsUokpWvEnqwzrSktLj7rC2CP5XHiqPlIWrHFuOchb2wMHgIS/OC8r/L8E2aoQZ
JfiT81sxhmge+MOH19JQ6uE+gJAhaL3TjfHGduVtgNCVozQZFrkZ96f8SkcaXCm9
nx/mygd/JqkrT6COVhaDNQgkCUQM9eLuE3ASscE2ujOk3U6ip78MYVTozNDHsECO
xGtYrLW873geaVC+DSd77W+Xrk38SywsZ991lnt7qdgH0Zi/zj+dO180VSPCvI1e
L0bCQqKMrpWk75oakA/Gg8/whxkagdgTWoSTBE+msPSycfM0eQ02wTx3meLTyXA3
sjOlIL1QNBThrbaXsR81aZaW0J3IvyRxWIb55xHgZOXAJ4KTuCRvuCRTc55w6J4V
xZp1P6W9oX0mq0LO8TeVlX+XT1MYnIZVpKIO6573LXeQjmkW0Is4BMmQd8pbRpit
0hsudprCff5rhnljenjTQL/eAVBzUBCg4mUwsLn9lHJCzE7Z6piiGjj5wBBBfFis
j6bKim1Llbp42AuO62jV+8Kn9c1yZyOULmA3XZatCLbbl0/kdKaErEQSW9z3AR5p
g4KoaEP+35xj0cJpExGaKFsutfFmix1SqKQydxsXhP8LlZmdjlqs7SBvlCF5ks6c
DqhfzLPMVbZAmasyOHxC2QxZEzDHQNEjBLeu/8N4TdXTmXIb26DhWrSbRtKzN14N
vQKxi3Vc6+iRXdVPhp2ax1o5Mfwq8aMzmMSnksHwxnmMR7V/eTS0DXv0P0yhmxt7
9rkN2GDyw2K8cEeKBJSgaOLqaN7c96Rcyljhts341r3J8AKF8qFmVyYuTxFx1ZMD
qyCk3fthOuwk7J8E+LohVVaPUTc4lon3iEruLmx/kKMa3kVzf9Pci1FNSIfKdD6T
Ta6+HnN/XHNz7+UITH09wgRsxBT/jEp0yD4G4UaSXwODh4B/wRne+1R7cA+6mhG4
2VfY36DZsvgCerH/uAuCT1eYNrwnaoHYcRq2wLfSU6o=
`protect END_PROTECTED
