`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Chwz8G+D7Bnhm5H30SpvzXLMSVRPoWPwq0MqNr8iN23QLBDTlO/KN13bPO8TUKap
UuYRJvfEPKTcz9bp9AX11yo9iLp+muwjTWgFdFqbI6a7UalrmKP00rsJQqySgdoM
TIRhh/QGOh0aS9wW+TJOKf8AOD+WgFL7EThrxvjxP4Zk42FqQbiP3hsKd1oGeTfh
zU/QwYU2/NCgHcs4lfB2/3cSXKecDEIMaaxbUIVmqDcMyjNX6lGCqdaNr39f2Azr
Gnynx48j4oKsb+A2SocsL4ZF+wDnWlfNhHOKIjJwGdNOGBHOQ6m/rkjQYrJtRxPZ
gokb/eWV5hnqlvnGXSRFgp7Cd+ThwNqywtw0FsoqnhAiWB6gQCt+u5mX9aXkGf7I
O7BgxnlhTURESeq7KaWJRaIpxWHAP7Ds/P29PqS/m0gGM3HfEaGUnE5lBiAR1S5q
vbz5U0olu/oIc+BbQflM6u9xTeUBC4Zi9VeTneODxN7YnQv1IVm1d+4DU+c/JB/P
0Kzw3Ovc8ZO0K9Q3hPgbINK+LN326Dij4akf2LaNLMWn2esptOjTbMqE5UmmcVbe
ZMTgnlBQbnbqK8bMCtDzDT71+FrWCzbOJuEz2XoWaDa0uw6a1XIiKrsiKkO6KWs8
eBEgjR4bYd5kPph0B/BlhYRkYNhcVE8B63Yv8eog0cBW45fpRwObhk3CYYTcOdSW
8aOuGr7UAJ26SsiXakq59XNcIzwSDp7nkPPshYLvDCWD+Y2OSv5TJY/GREpBKh/1
+sC10Nry+qigMrvutWfqgf6I0Ka//wrnMuNoYxiZjWJCsJDtDioio4tY1WPkwawE
6QOaPkuumxwrM+/M+m23rv9uVjuuT2/3NHS3VimBRfZNgOmXp69hnnbAN3sidfuU
pStPaDFBHWClh0zWbfeVZA2yGCuBlWG+YK9MQ/AoAQvANTbmUv5s0ZIIrVIEmYQJ
hofR9qg05DzNSeE3blQrQI+Zt0h5DKO0lwe8yukLqYvBN0BjEAWP1f7D0XuhqJjl
HO5ZR2PsnBe2hf3KkEz56AYFPJep1qgkRO9nA3lvB8Pyz8BIuonuIII4V+hIMGKa
Tw9UlagGBFvvD17QFuFdi1mBmxULI9Pl5QpCm4c3CUTBDJxUCsnxvLomDeOdmtAg
utwPccSC6mVrqb4Hq2muKND01XuBWnAIVVAqoktpMieEjrtODxVgIUIydEOuNyqz
qvTx4wskPa2a+TTV9lXZJCdXVqKOetLqQrHNMhWdqQP4Z2flc2hEzG3HhMR1yXnd
ktbO7jnqmYWuN0uQbKhIqiS6e4MN4NeHaoSC86t7wlcebMOC8tLBnyN64zREKcLR
VuASphYLrfT/XT0BhNExnGHF3hSCNzASUhcdLigF7Whp/lUmZDY0OdiYUHrmkdtb
izX9yEpP+gsrm5R08mwrHLpdx8SMF3gI6ITlRx3wh1JdWGAuopstjFxyielERnEc
B2li2UGZZfRwDpYp4ah0MQ7kCwaASmwc3PU25cMr5Er/FJQbN33wwOSVuqmoWOeb
wuRAJKI9iECJO+cCt9p+ooIoxOvj9LGTe/gTFMpMw6foCnoS5B6Bn7hZqdbi4jLV
Jg7i3a2bR0hAkc1gbFE4yfMXnwYdmIL72jcz3sq9yYzTmBcQnnLt8rss+u1xByLm
ZVlBpKGiEc2TC67awz85nn7HdvVbTVIrlpgNO0XxGz/F67bRxlcvYj3AVC4+zI0q
n+Iiyln1Vd4U5AlRUm1v7ibednpulJb9DBSWF8JbjVm8vPcxMcPVSe74q+Dq67Zu
SGHqyMgAe30ab+ZS78dkS80Djk/sIqiZz4fA0fbeasYKI9B+llYOZcV4qHvfSjOf
PVIdx/7KdxtzljeZW/Hi7F2uxOKblvSV5/bPrjLBGQMgyBDLjLT9OP1+VNFcsCrj
souCe5gVEYetYc+oUgQjKK34kTEtf7O9gviZH64cvMFpVgr2d7IfbfCCKV1mMEE5
1DRXR111TXolF0Nf4LR3IAcRdTCTSvZiv8F4cAk658+G6weXfF7j0bFIZyhkN3JL
mjj9Fae3z+cpbEm+te6vE2B8ZNnI7rqIQHnLjc0w6BAMjfq8Ex3v0XiwEZWQFdzm
De4klklDG5pvndbuU8OEwj9wgGSevP4jGBRv43xV7oi2tftimFVI7JDsrYgyYKpq
DH1BjeEYZhXvZVqg5KZYYWg4oovaZLg2S/zNb2Q/P4Vd3Bp/Pg1X3DbKGj9q7rev
MiOIticAbDwyWb88gqn4QC/YhhSuiptW0zP1n3d9FOYiE8Zt1Gs+7Fvv5hWQ+on/
ojoXhfHTOeitgx4Di/IFDaOQJG6rH2NPHBKWt+SrrPVJ6fGbnLjdCufGoNN5ZL6o
RHYcj5yEj2gHaRNru53T9TyIol5OvIjNXEq/ext6UJ2QgPJt23BhFSy95aj9KX8h
fq+iTefwjtpLikJ1ESss5zjGhkMOiLjZANQ/kGMT/pvU0gi2AyBrdG2zqpmv7SKB
6v0UK0Ji0VfNMxI9kLB5PQ9FVWMrfVDW9BWXdWH7FBLU/4R3dcUv8aSsWbFsLLyV
cUFJKEaGxqieWU30Qll+DnxeLFmUJjocyp6oFpMlOU9xCIE1L0wbtYmcHWgRlMvR
+N0CtDA/WtKjRn/rDblBJiCNju4Ay/dmbZaXPhZzhuCH+i+suFB2RHheueZhIYDQ
ojjMRUgH0XsGFJxif7TNiIWz3V3p0OlIO41ZLD5W5HaB39RRYgFD4Z0Ut3B2HosK
9jvh/lQ201qtPFXxhlXdGkDSXwTpznLZfLqBCJfb8BSRGfQpp54R2b5Hw9G6p1sw
RSDzkVCtCTTYpVzYpYlA/sPKxmnbwPSYdS2BJEOmsbZx6vJIc/6hY4NYuOG6iqti
M36rqWwbAa36xyocYcZzaDEQeqGptsPz2yhEHtbjgfnSzG5AyJLVz4nWKUQrLjqb
zsc9zw7rFKa1J9+iQV3tenecqlnYL+Tv64KitzT6zxofpm5xAs4nx762M6Wfe6aT
eW42d0DXKzQ8VezC0KeEXRyeO1EnCUo91v91CH4DIk6U1lThcJwH3GYnfJRBfx96
ZaqQd18NyYcypC8Om8hH1TwNFeN6a8FjLlAlgXa1lSvKdDTHmHcAfFrWYmoIQlrE
nQb15tcLkUMv4BtxvkHQxwLadbsVg3isbXiA4e4o3gWge2s3O0/97gYjeiv+jZO4
q9xHrLHUqJJfGSwWN4udNe6745BZqtQ1qnAShonxez+fzIXf/+o8d3Ipuum/5D5r
9fyb8hqCy+iYuYTfGpUkCjftLmb+CoqSFab3F40F7TqU/PrQU7f1Mg/vBWjdqzYO
fc266RvZSzDExYY7nG/oQG4QkXMlZmfte2cnbQfIDzruKareAjDUCN/Yg7vIs86a
gv7AZm0O4qjrfTn5UFtwEg1BbgS4EBGk3XvR2ekINQGYWykKbRYV4s9PtcT+qdJd
3mLMiaAdm5frsu2fjHku3X7jBnhtw/ReLwCfbKItHx5WyFzuMzE/GEEz2G7Jekpx
OD54AvO5qOJR9BriiRF8RcwpcRlqqQ8NRYUIJoMGGTPCvwUIvxSbp5GAEO5qT/tm
uYTQ9MLUSjd3iUCuy2kxhaBV97bofPHixgCYOeWgRY4ehtA1XIYYfeVJLcEPeIKf
6KFlzUzRj7ipgn892Pin9H/A+kXpkGq3HgJlzh6r0sRqVI4UQF8Q5d3KkrPjfYJu
fmQldAeK1gPG08xZJ7dnnYFrSAPP7rbQVjZQA/XyBAZJWT/TasT7egrQ7ScD4pAp
qHrLVM2bka239J35PMWu47nBOQ3kLkrNoPnM3KC/7go61Ii5PMS2DXL9meaWEboW
9HaLVITwSzwNxlVZkqgfr481p+98LToQSc4eQXn+GhZNYhI4R1iW99BhbVB9IK+S
miLNT25ST3stwp0BKHHTEH0n6kWU4Ul55JWuubf+GQv5RZZuERcQLcJ3sWD93pO0
iXkO1tutHeOcVWf5PsUGKTBeNDAGCtyYOGF+9rL31+JSrGEyDtJuD1sij6T5NNkT
RHU8pPeyoHR1sSr1MImx4Ye0QAhrTnicI8K2lbJQmV/8eFnPDJGyTpL6jEyZAEpv
5ssBI81qUZIDV7gGzvjiGnbODU7MJ5jmkTeNcEehHTvQTP1UlKc3RwmI3lgXphPs
N+MUhHhTIshjjMKLu/Ye+gDE9hvGPNcyU72Os10ZU0kt62hsNqAJ1taRHYhNLY1V
NpO/h/OmQDtaO3jutKoJmORBXdUriF8lbrmlSq1py9GvUg+MroLm3JM8wJYUppCa
4YvTTU205G9h+PMHFQWkleBPIQyT79T5LBSRHQm3jh7OWBY3O5dYhFoTlwORssUc
9NaLPk+Wnz4mhByeIwEwQPjyJX5EiXvtGSvF+oIGrft0TaAZuXCFct4CRYhrdfSu
taKWAe5cXwxdG6bFexLwWyFeEQxDXWxvXNzurb6nipacyAf32fruEvzyyi0nH3o0
kQjC4/W8VRAIxmXYPjalOnt2oC+GpfJUoAloMAT18qEvw1Sh8lUGdgmv+JjH42UG
1W00q/QaC0/ARf4M//lSKhLwOIGlb0sgU0zCyuR15DiurSNOT0WW11asw8wAJDZC
uDaDqIEgBO8Y8RQ6X5QGzYSjSpjOxzDJ9Lh1rms4y29M5URY/Hv+Bl6fftBhzrhn
w+iYsFJwA7S0ltC/wm6TrYYSH/9u5t/I+mJM0/zbGTOqQrFvcKHddc1NYqprA7y5
/Z+IetVp7Gzy8mZ/dW/AdkIHF38Z+OygIP4j0bp7H1uDFS4pKUjpPqdFmg+UGBiy
Hy2au/UpRmyAwAX8E0vDYx1NiRU7YIUNTu8id02+47wfOiu9FvIh3tp0yaJ69ZMn
jQ5LbdlGPDkrLdwMVi5oqSDmLUjYIo2WTOUZ229ZC9QkDHnrHdA+ddhQDIdKQeve
vzoOEPLEoG2PY76L9ddoXRd8HQapQdeDJzzGcl4LnyPrhmQz5j9aa5gav7ZJ4DVv
0VZgstosn9YFibElUBJ+aSF2dGSPoF8ARU64opSDas7GMAKX+72dfN8NfAq4N2jP
MciT7VZ+G/Wxnr7/Ev59OHFLu+74mJkqE4Ub8EXshOMsRcoPZL6teowH8m+oBJmS
L9Y5PUFeNiDrbkLVHV57XXnVd6xgQCAg+8Nlwi+5ZS9jnlda5D+XjwW+iPtS/i9C
1s1hcI6uXjbClL/WZebZnhbEaKqbHHyUIfUTps76tHS/U/XtVbtbSInCvPElhW+w
Mk8hCPyOq1we8h5bv43v548y5NZgdTA9Lud/qCYrmWTS8n7N7XbYK4bnPdN7CBfx
DYRzYk1A7ZBZk6752nJzkftx1l6IVsSETEr8Lkmk23xYzWioHgVYPZIfCV82nLZC
7wtSwfesAwjUpF4s7ZBTD5XMMk4UmsMQFPgKCNzdRU5nD/nP4s4dNVCu3DyjNNfI
U73NxAgTnm9G84bWbtjwv51NvHhpteu4gYrM4RiORzSA129roCycrlkGBI1Y47fO
Gpp220fyhqSJsgjjaz6zzTnPqBfZkWA1DHh02V3hbdFjEcl/B2iej6f++iha+t0u
V9p4mVFBVCPfzwjWWJNB1KaaK3yvY+35GfVLPnckf1kxidhJjmA463nFR8M4owJw
YYViGPLzuwRhzsUemK8+q9PmTbb3i7f//L5cw6uf7DEi2FosUsY1Ef3fO9IjRWuR
xuz2uzOo41mFPvDSFptlS6YFUwVnFKiGObdmWTyAiFf1d6mCGJg5KPXLuKkMyFZz
J/xrfMkwGzwjARtDpkq9v1rHDVBtViJ8bdhjJ3rXEinkUTisdLhpQs2zmilllJVa
AcKPTGVF+nOfJ9+vNP65WWmkyYrUF1G/UFB76kSh8XB5dptG4xquEWMCtbluoybC
jtpYQ6sfjjJX/BAYfSDZZ4Hs63V4Yz+/OpCxC9UT2SmTBgAAUmerFMjQUNs7ZmIM
BpMKBBFiyc4K2w2aLKLH+iypBp9LY0rt38me0c0AbkO2CMt8o6kLfWUkpqOhntQV
QxPO/VOzKj5JV+erPHjtO1sNi/ExDo0gEibttOjTHk0=
`protect END_PROTECTED
