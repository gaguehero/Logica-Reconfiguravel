`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DxyjqbaxR66k2knAh0ghqHRpwcU0n3wl8p9DjmKEDagLzFK9tH0tZFDO6Cz/Qnq
qovj6lBgXlisDchw80X8KcdSvzghJLtmzNK4YVT4l6ddzhx+4AszFmhre6+rIzTM
PKYPBaO2EHXWA7ddKlepSF6O5QLAZkm3W9LEsT06Xlwd2mF8tV/XNT38s5CjJwFs
+qcyQaTFin6O6kOqxEYq3JY1vdDlNi+wQNoL/K6jhLw1F1MYjJFwKhevbTMRCZMv
CSLI1fJ1qubl58M+b5Mmy8rVCLDhYQpivuAS77f5zYTxhTO9MF8PJxbZal/zVMAo
nl68ix0+ctILgceOdcv+ZdfNxDSGXxuxcuox+9wtNKOTuwbbmuQv4132DiPLj490
ofxS4Y3Lk4dzMPzjxVaCxLleWXmPEgqQKBFFl79ARuU9SToUez2eg4VZwiOVrja3
L4VO16CKjLLDrgAwymy2BuSTRzqS+6+IxUcZYAwZRN02QcBt/NZsovsoHONAhAN0
XlSM6O3U2D8RsK/YdYjiFNb1d37pClAjIK30ogQq5wPlDMAtdrF8vGaXJmg+Cn37
J9hYq6ZqiFacAKVVIkvDA3zOefwFbv7ZVGZivRmA7sncc/88bEuwbBj86/8oIAcs
Rtxw5f/sWA1NFa20c9v6AFgwrlBh58XG3tGd5erLrBNKwXLA0pMWg2rPiQSKQHXE
QlE1ZWVKOEyXAaKV0rr2XJXTfeAP0AGQD5X3j75NyJre3gbzpJ0LRMDyRP8nOSNc
QkbGa7iOudT15Iank9XdalKiUZ+23vcLEP72sqLq/GAaBkvk5fV5vvNfItlnqI27
RtlZOH820P9Edag8O68Pk+VGHULthrMLe6EImiPvGeQvFfcfZunTM7yw7akL2FHD
6m/129XPDlPvjQhwA7IukRT5CHRXlnMMwYxpUsnCXCMe+MJ03cQVNiDtazOA3vMd
yhTV0n3aVdgRLTvxUugujx4IieBdeSKyr+85PbdiApx7ZL5sVVqeBGrpf+8cFFSo
IbT7xQ9t91H6keII0W7qJhhDzbho7Czmlc5dqCvhXQgnNxrJ6CnfyrHZaATvrrN8
E5zbllqoOuwyFyCbqp2j3l5wz1iEHWKOzEAvzLGFCBLD5hvvini0Q7BMth2b4Jqu
fZawTvy9n9LobnrA/neZqsqpQZKALMytO1b1cvYzN17ZSLoVKuWroE3WKc19k15f
UkT0aqXstyKAjfz0jRq1NoJPPd0a0jPr8IbQXfZxDhJMON2yUXONzC9K9KeasVUM
E731ixdyssdf2qevCRCQHCsStQo36THybFJYCac5X0NEwiAbV0xtq1KSzGY0tum4
hnloL1pZbJlgTBHJhQO22O/pTsGPOvbvVLLtr1ssgDORIusBNDwZTQ9qhv1DtLjX
kTZ399I546XSwBLeiN1KuFOIDu6nzfQG0jliWpbymXrcRFFtPsavLasPBnVW9K3u
DaIkytwmnF8CkHI13G49Jc7eHwRpbPt4Rop1/uidw37nkQc+1aFenf48ax3VDB93
sI0J3Fw3ZlUA/seSooxdPZabvRbnZfVRegLiTs0g6ABlLSFy/4sbLRpsQ6PJrPLl
2w3r/givSvzLaMUBgdkiycXzocwZWC0b65xVmanguCFXOjWHVLBuh37FMmtADjgp
jvS35Yj/U5SZuq1OlsEfg0iXDagwuWj0aUceeqaZh3CRLbxkmPjH51YW7XoeCsYz
fijVCq7UidoPej9CJtf3zUZPDfLZWrA+8LEfaVsRJQW96Zta0GSXT+VdLZn0UeCO
3Aqh4Qf3c6FvWdj2yH6pGVxX5MeAYPijSV44SnJIgrB5k2d0jGIaAuJqLpMbIx7Z
6fENUVM55d4Plw13yamn/nlDqenlGdXoE6Vjc0Onw3xBPdWHMpBBMmlUX+ZRHLQA
PWf2LgwTr+H+g6UREHWl8sPfBUH6TM1ljRxUWnVT78BqrFBrWh6Bh9nVNbkoHjOH
MixekCMRl2CvtPPXwZkNjnUyRAOAGeOVUJg6aT6x0ZRwDIRAXM/HSziE4YY3PYRJ
ODhfbRQOehCaLaQRPTJZRhdFTfWaeA1o5ecRSff/S6fx/bTxzlewAIhQ+A6UDUR+
6MHZ54N05Try30S1yq+W9vU7W1ZZ+K3PBHzjFDUXsojstD887sDD0hW2fTPnAbS2
Fr6G5KDDb+WEAChdy0MJe7mrpNNnBL9QDTI4qxOrU91Ik0FJtpS+xJRMBBlZAi1m
M4wD5o9hTXuehwW6XNqmnA==
`protect END_PROTECTED
