`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8nl1KEGPP96ytnwqubGvjYYvfOhcPATyBEn5hATdZdQiGBYx5w7OgZcERRinsmc
a6rV0o2g/aJMh67Gs6B5cBFlvrmhuFZ+FTZuk+Mfsw3W9aBGHi0kaLvU1SI8w3zZ
YGBMkcVLd21uBWKm1jXIWznGrzgQubhY8PsuG64tyVhSz1mpphOAx6WPx46ELL+6
MRYQB4Nh+6LCCWjrydIHUvNSJVCKgK2+Pj3dZExVNdJ1FQAUtgFD+kezLjf6clSY
krIP33Swqg2auwiPhQacF5TnFw+ZkVb8aBiacCvbaffKaWq+6ONvh7Z/D+XlXaYf
/W33Js2+iqYCfCCbajgIX5upLLuSI9gfxcLSgNZMM4aoboJSma+9DJIAY8fNlDVy
Pny/ooG3fx/MvsYsWYzfy2DG3Evmy5fEfIAEzmK2NqqZpj+Pil3UQzGFoTIonF3f
OeFLXRFzQadGdpYwCjhuyfi0MNAioa+gQW9+jmr6yTU9pj6C19zobCCKBncRtCUI
TakcPfzTLhG6EeSUa1TOo/U3FN9ssCIaglddQkUueczf1AmXsGCd0mqmSf+1yWWX
NbNse/XI5KYYYVC1YAVy29NpvkJ6JIsQOhYkiH+L9NIlcXpSFh+z/hTtrg/AttX3
oJoJGJ1lsAzyZ7OuEzG2q68Ai5A8ubFqC+GRRxAKr1e+dNmnU0hfBbpQPoyNVJxX
W74EUTDHLw/QqT2WNkihnDILQM0vjUn2XPHMI7Jjz7aYFRMbZ/C7XwA8kjvkl1AM
OMkf2Np+AoV17B7HXjxFJvXu3KEPVPMp0H+mAiO+21bdvuh2AN+/UJJSQlIqgzv3
T/YUMNXNHoQ7gBpvqOdRpcrIpPM85YJHZ41GN7/xYP9VhGGa5RF7mY0Oe9mMEewc
rPXRV+wB8/vRK8ORs5aYicDtRsvpXXY3l3AwiPEDLwTO0OPBrpuceY/mzqDylKLk
5Oc3VnrIUMjljYKgphc/2TdAx8wvWn3BgR6/VvFJkpr9Rll5PxOzCcVDhz/vQp+j
jjyFO6Kh30TCSj9TLXDBSNv2EUNrgagE+wYkiCpasYzLvE4P7yZU9Yu7AZjRt+KJ
Jnehydpa/2qxucH98J3WEScSqdW+IscU0BId2fhnLCpMyP+JM+XQ3tDNNATT8PbC
Q0R3VOZuSVpJrueQRxUWPM15M0L2W/2cmB3cZ/ryg5uvTuQlgtEBMXWZ8v5G5SvJ
FyUkC9FZ1tX6Mean2OhBm98NHE/H7u5/6Rmvqb9FPko4m+yMXgQSSbdOUM+FafIz
J8CDSaXqIrdiu68Glxsb2fqs4QNannhlMj4YFllD2vBWMXdKc//EHzsM7YtPR6lz
ZfqjfFAzr7IeNI+hwuAQ9cUieCC2JWPAjw/ltfbLaGtloHpqzb6/ijVIwVuPjRT4
+qYsovyqT5u9Q1aGCCCeSGA3Crjsob0XqzKEwPmUSvuUczdQ9GpHyCaz1bCImV0h
o1GlBwTWn7Y56oKBIG6JohBHTy/ZaZn8ieC/HWOIFbiOfp9wouep4+7n9a+SVcwE
Xv9lDUXCaduLEoh5L9yjBd+zS4lJmc2toKto7xyoZt7/EgIevrqQ7AqUOBcwMKsy
8XPvTOsZruxTJJZQzaZQB2pz+H/qi49qdZj4RIO4L9uK+tvH3AehSAH5mmpiYOMf
J2jEv92eBE2Cik3xYJC+q5NxMb1HbTPsXjPVJ9B8CPYjYik9tdGphpwQxIRQqd1U
CsPk4q4sS/9Co05/wvtxqM4xHQk2bshiXMUZYqabcFt/cDLTzkMIdxUruTFcMda7
wvPLqxoYvbMcR/4IpIeQXqhOQZdWx2OUtDvsM1qum+ZYJLlZxlOq7PXhdJFRNraI
b5GSjbPMl7JqlaemjjJeuH2/8b8EZOwV03kmugxcSQXITnLW3c4B9tgSCYL45YXl
y1jNTWZCHf81nS4UlPPxBMTBvP2NPoOmKaEQ4ETcoqPv8tpax96q2p+0ss7Gvdvy
2+2JJFBQIb3eaZlvIFlBAyQDnY/UeHdy2uRCylJAUDnVdm/l6CGrEKRtdq9tA4O8
QtoVjyAYb9dIgG4g8tInBPd3yLYts17Ez+WnzKvmfdBhAaZ/AHmiH5yFjKEyZRq9
WoUVBoljtpc0xqzdh46TYJjaj+swAgZ0uriB6pN/d/BpxEFYymXnJ07Meo86A8lG
aaoChJJb6MKs0A/Z8VBgfS/ZiKeleoKeNvgVSly80cNK4ZILmL8R3gICcLi/ljeD
ciTwpJ+RTYgzESx0YmD4GiBEPoFPAfZbhVKe/7DiVJwSIC7mEnDsVD4jBgbKYLL+
VKd9jYOFHB0tRMeKzki4J48gqfJuWgozS3K9SjtT0l5FzIEEat6qKNyEVeLdpVci
Lp161Gdg54KWICRCYiApvflsTbbbhT+Fd/6N+oYl4VDZaqp/uxwAA9TPiScXC2vJ
N086O6Mx7Gp3m5ZBQO4YO9xn2FDSysmJpCQpEdiytZeSm2bgJ2mxlG3dg9WjqWxP
SNlQDLE52g6zDxReCYtEJwEonHUb/r0Iim4yIz3jMqCgCGWBwuJJ6QJDoiHYXHqo
hmXrRLqj6K3rQYT1scxaoUWy0L40ks5i57MrubDBbkNZAXOj5/LmpEzx+toaeKMl
KfOfcGQ6I79/scp6kvt0kfwK7WrsCAAWOAKeHRXOxov0MsCzuQRkSbgOFCJyNw7v
1/w8r+yAN5sDiK6MnOaFM/KZ0wA4jH6rRoX99Ea+LMjympmkUO815wlqDeGPbChh
BXb69ivqY70e5jFF1oaP0mbgEaq3iDKMujFvEij7A4M9TBDhFwJ3QR4eOPgYdBXO
f18GLSqHnZ45PcQAO9XQW6w4S1wkBqx/QMfZBrZ2TGJnyx6yW+OgH1ve8xTQ2sed
CUw9/YSv4bYEGYfHL8+YDBT4vBeqWCfZh4o99VGh2g8QMGACgl37Y5ozcPXDzmGM
zlkz9lTWVucSV0U6hUERJyRWTGCBTJWYniujlERrXhSJHp9nxHYAWPX/CFB9cANu
wmsp2BgX7K/1kTeqh7Zt+b9H9eXfrtlp9YG9KUTy2djmCg1MHVBJbewwkyIPdn/v
Osp2GlPuO5ImyZFZYamsUDaiTAGAW2lATlmnYvP/aibwMMrL1sNF9ggzDRVLS6KZ
mI4vNh5jka7rA0WdXx+0xpAc88u448UsWO0FslilMGTeuJJqONFfCD3cyeaFRVS3
xkWGaIxQp3f/upzQIN/cuyqc1rLMYW9+734rsmSWTrXHRSRBQmOrSauajmFC+y+m
lKSSiUHU24i8DuH60JPeNcWDp8kKhqmXGkV/bnAQ+UAqQFQKGIwi3AIGt96KfjkT
4uibLyJjkcfp0XfiPtqBg1BDHHGakNObUd5zClvqzMgvq2q6wOKunO6MWtB0Ajgp
JSspCU6Y7Imi4wSLBjJkYtIC4T3a8xExGLUxs33c6y9SuBTD2iY4UoHexf9W7S5R
0C8rldicZ5TlXlgCFyL+h68hFHhsNlVY+ylgd0IU236zT5nQvFwSKXnVJquOi34y
tvsXm3sfHjogrDmI9n3bGB3AdPJhx1weZPRO/cjCTviM585ByfO9YwcBdkQFKKoz
zUDR8TzC7Y+UJGQz4hp77heqKflXAYfcarlAKkdK3T3y39twKmqJbbsiK8DVjfon
nVA+83vqqs1abnD6nHQ51tOgRAWfAKCRlyaTgT4uUGd3oo9hD59GcCfv7A6s9jfp
sbh+rp8Hk9WfIoz5uojPKTIKJvKT0Q+mxNdi8mdFjM9MS9jFydpNtNzUxde1jSKt
m/pwoyYUrxc/tk2g2cttLDFcwh5EqhWC9fk+AZjRj9s0WaZ3tCzOD1CMdpH/dduK
sbQ6mUyJ8GzKuwYe5PawsVEgwEUCvBI5skmzoy+uuh6dZ2q5I7BO2rfMFL9hzjp2
djxm+wFiqkcWpflIYOOBxDm6H/7yAZBsR+621W4gibVw8hkvqEGWCjm9V4G5uynZ
aGd757N8pa+0roLUldQo373ibCa/6y5yxaMiI1S+hQT17dmL+HVffpsBZebTobv+
aEt4xEZ2h0fcbUx3g6oiXVewrYuRPBIJRWzsxpgQ2xobDbucGpfraH2FojyFPFCn
NKUuDTwMFEIbdysNEYFifdmKPx3qFMd117ybG1JyZWTkoRWgEbT44Zzi1CpZfNWb
x6U4EUHoKtAKOVSgHH6ba8TlokMnuNOyaOxGPcUKZirXgqcC5/ZP+2gtH/ceyr8w
MAskNi613c1xFj+3cczJ5t0CFv7xzqW8V8GvAZgFga9hIuZR2WFM1EgjTPpwpkRk
amm5zNvl6b3sJMed5AvCYz8c9kr0LAqwRormyy4p7HWI82ryM/kfBjfi2LoLdb+k
ZbETrDC1W1YyGSgkRUGyol0t/161PpTKqgrmiG66bnL8PHOU78dspMpj6RzMFIzb
GcXmfIgvQbcxUOxOnZgHBhWEdvSEeSlAoUfVL6X8H4YMViXwchkhQ0pXg/s+NK+X
EPedshvGLwhnlUKbRONtNTH9/LhTBbldv9rPFTHvXq9NG2iAyRb5qgYFoPLNp8/U
mQ2bEyvXYShBiWyrL0iiSTD3VyedbZfsDUhnYqdo/DeNhXLXcHcubzaFUKnj6axa
BNFJU6YD40qyBXo7IGWfndG1e/eIWDWWoB6+46X6pTGeqnfOIE0k2KP4bL0dsy76
J/IFtSUSPQqli3Ynx0oG6imvAvdo9gHCxrtwXgMy8RFTnfBWYPGMoZcF/M9Ic9xl
H34l9PPEQRKopecCl6IXFKwTUwmm+8w0+FgpZGFI3QypSgBJP47mPDf/aObGn30A
tirbjHDqxmg7CUA6FWqUN7hWn+zFgb+GwyK9slVpPEieWTjqzr0relSMz0d10ht3
6pLcJdDzFacaiyzuVVH/dviIZHVbeMt1zGVeLGnADiduIZ+aHIG6vU5kNQs0H5hP
3MwCTh/XkBjKnZB1NErBd/GsGSApT8IGAzzkJ125XQOeLDx/8WjFaQ1fUALN9yym
beAHLhUMHBl9Ic8wk4G1lMtSR3zoyjb9YEYnp7r7WpNrmmcwCkXv2ZWFLSpBeRiz
9CsX3++wXnjChp/0Xo2R3Cj2UNPjnAHY62Hd1jWf+7Zu3WvvKVHIPTNrSm4OgidW
p55OfQ9qxEisTvFxCiGjueO3flgueT/87s+/uMhhtV7PtigbUEaUYZMBzsoDbMv0
rlP1rBqeqsvBIZwTywEP22IOFmkujYDZDYxlycH6tqB2moMkY2rSxQLMKSm2hNn4
/BWfCUgDg+KCJV5kFiqg8pSXX35ebTWj4EY5GP5eeFoNczMKQM96zIwGjwfhl6Lr
5k5wAOySbfp1rWzwqoEAYf2udA2LXxkOXVxyRFwnAEuFaPoSvkA7m9fSMUXAEnbj
X7fqIX3jaw8s+UkdNkdsQ5SXk5zY6xYK6IXSmhEVy3469BkYjkKjj8rHAu2A8lMt
QbAX1TXv/c5PfLRHXQET4o52lSvB7XMB/Eb0YWw1ZC7GM9uo5or0YVSThZ1gtGwF
GqbqrLCMxrypWyxwnf0bHrb2z6MGmF6M5UZJbKUse5kI+124t+7nZ2rqHUOqKHGJ
9a17EbG0zfEREsTqlTE+NV3S++ONvrSMZYZplI7GkS91oQh2zWtVBmb04VXIb4I0
W5sRRMayo3a+XpDS0e/ilfAwrIykEGLhvxuRBvmZGZ6kNLBZJvq4T8+p6EF0NhIR
`protect END_PROTECTED
