`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yrDQ2xUpNyGje8WoE5Y8LczGL5++S2fhKiYcJ7sm0geZrNzS4V7PjQL3R0APtQgH
erJAlWh8CDL4x65oscrrq0PWDuwuD852DJGBoTagVxqvxzmgRKcR+4KX5VDF3Jf1
TmsZao1PK+25JTTsOLJZTGkfKTEThF9Isbz5mB72dWx22bI80lCqwOIpyuBuRBZL
4+V/nLqKX1e0ntABhrAhIqsRF2YbUgLGz0QD3kkgl6iyAJUF1b6H5cZdD1iv3IsR
76rxSKN4yXpOg/JZFTxa4aN1hNN6oAtZw3kWq68W9JYwttZUUtbhMK43C58za8uc
QHrgG3VUAvMCJEk0O3ZGBNuE7DUsH42LK1yvQZJktvE8nErwTrsSBjyOAmPc5ydj
hwJL5mWx4hhd6CUVfS5tx8EVlW/dE877bfMygjnxHU+7F4sGFCmJNVW58jeepZXZ
8Iz3qA//8BP/CeMyjwzJEtDKN/XR5X/1YhGB1SyWFVN6FWzJmhbnzV08tOR+GTpl
jzAPQch4itJzxMuViZtIrElF/Kseg0TgTiegnRQtwzuCR8vMbRyJevAET2E2iN0U
aoo1au0JAtfapoHsON16FYamPwfwV4AYp5r6waDJNI1tlsADljdrgctyx/nVUq6E
emUzFLt6Vu/M0/ia1nm1V9RBXTvS9OfLjH4gakLxf2kAlL7gfBBSq3JlPLwRQMto
oURgIlGdJ0LaxAcxmGJ/j7IFPZ6aMctLRJcedpvJsal7ZPfvVnv4QRP9reTo3aOG
/2Z/YCcXLEK4csvrg4N1PVunZ8wX/ZDRv6SQ6nGZyHmXGIuIVsLeuIO0aPsyBglF
wJnqbf4e5syC08SwZu5b1vwSGHfPL5QpAWwEZMncVAGAOy+R2EBFBeEGy16/d8zi
nEIcycpJVprxRTmdQqkOqRSA1ax09Ssm26sfilX+xAicbl4q+IQVGbg3FWPqY4m0
dWrmleh//vvIBp6XDdfajO6/kfQd9iQySgC2BWxDRBqz5Vk/YRni+FiGRnWNNtfI
xp19U2IYAuSyWFDg8JpzYjB9yoooLRzzg+PN175GXRD/jVFdUvSjOhk6ZMI9LR69
Fxta3WkmKvem6o+gNqJIQJ1l2lD7axwUhwIYsQKnnlcQDke44UVvpv4XtJa8dRFx
Zm1sqhpOc1i4PUmVmie/yHyODVRdenerwIq+P+UGCASBHoByMUslFajmRqiMQn1y
5AeS74xcLYwcZs/E/pWLh0WziBMcODhwZi0WdBbNYwal+CJjGMW74gq9u8/OI4TW
zL8/81IpXj359SfdozjSpTFV+XPAIC8qoybm4T6UVAjF2s+cC3wAMgons3mK9h46
PKK2s9mGwVSkS9mT2PGCeDziLeE2RIPJhOW3KfJ7WicEaw6gOaCKoXpzlrEu2PH3
PIyUr82fN0mBIKsX1f8vw6xrcC39cCHz3EGrjtImIi+durnk8nRf0x8y0Tso9sT5
IiCjd+6mjCUDQCPf+ZbVeYrmXdtu17s2RiYpzPhwfb8bID18PXGsLhkS/0paMvUr
/Jd7XNueiyqNtdPWRxhjOi52dBjQuEHSXSsbKU8EbXFbgG+bgK4SKrjfkNM8JH13
qF/xmqVqSWlqeJez8BsUWWPcgH9Pi50IO0Xbb7m46yBLjZ64MM5C03M4mym/HZzR
seO4qi0tcOdIKEC4p4HuLaNK/CAbUbJLjmceb1j7x9trm7wa5U/aqHp2NWZj7xZ0
vRwevjCDTWSQLhhiHNDuO2yv4rX+xA/UYIVpvzWVnsc9aXat1HqGEH92J+5LHvSn
UwsN5XtjTrNJ2ER5O5HCYrl8/7RSuaR0w+7hVvIQ4G8NQXBua4Tin90jcDWZVTpl
q8BEoBVToKT78emh5yFuIWdim/eDGA15YP/zKLAhExof5DstKantmWoWh/Vkn05y
Ik+yI5CkS5vXc1WdvLMppYkF//x8lKTKv0qEj9faXuVB9QWAZh1zfPHi8RIF++1+
xGA2vqnov0EfMS9R+EWR3qM2HLMEmCZLfH8a1o6bpNBVDaigTNd7u7n96mXReQ33
7P0CBkpRKp8prQNJ5FDZSGj+2WO837WqMcqvSgg9ARzfMrC22HB0mb3JSYoAst20
/Mv88+UjcXm4MGkFG1gt9f7N6Q+vFQVzCQgQSga6Ara09pe4ivvmGOHd0N+M4QvB
R87lNSdRFOvGXJ7tgnuLaDveG2pHQI5ihwTmWZGo/QVyiL/b0AoBxN0EGk+z63EO
IpSerQ2gLp0gQ3gvS3duNqUhrvsi5oI/S5JMIfqX2YURB7yT6bDAu2mSBaCEUMAi
LO3wtOKDNFHk1/7ccxQwF8bLYKKPBr8brHR2JCHNut++Qq91BkaPe3lPJBivEPrB
bqsJdP0KeI5YRszXg7eaVQCz1aIFRNKk3hRlqU/Va2VyTHaURqCLhTSQBcQFphbd
teRq2m0JPbQ3zAS7wr7VlpvuwLmsOovWXlHDaJSgLZCE9Cs1oHTPFOdW3i4+bZDo
ZBUs24ZCfW5FY0Vjm/XjqloBuVOO4qXuk939iX8mFzZWZHyfyB5gBLEw0uof01yE
BG1ObCOT5Dq+w6P0BrzlQX0if5LiBUh6exTASSWxIMLiNHQTRVV+O8rPGygZA/g+
biJTChEBoCu9KbL6hXq2iMHRcPwSyLzMyDKGfaFsnH879DEjyptUhMQR/V0pvlq3
okUo6fBfUDKC8I9dsnU0GUqUE8n0SLQx/iJEPC92cgRmx+b6il4ZK4XxIXajUDvd
8qaAGPx3zditvBIRTWlb9WsWRc2tM7KqNru56FO2uJVix0Md9LOtPBnVAMh5Is+s
HZjzuVLhzDyZBuQ3b62KIBgjcfeeR3p95fgIne93stu3WmFsCDVLwbBHUkQ0RIIA
P5ESI/gnQURI12D+pvnk7JrEG0ukLgGYk6qMpmdYylS+DRJwgMiSHAbMtMNTKrN+
S8tYQYjGTOvVLzhWyglDxRcWpcoODBDY1T1VUnXOaAjJMtJe+McXTLkCh9vv71YO
IKy8JfWBXDOq9mUVa/sY3/t6DusKdxSKV+m6FFmOHcf7ig9tewQhnKjLyIuIeuN9
swLGbGtdkefOwEGUguhnLhfo6JY+Lz1+cmHAGEUXNWmoQU8RdNpaZOA3kBTeJkYM
uVqc1lV4ql4s3Kn0vvz/1FvlcAQ3RtcdwUZaV/YVceup5xJGKD97K8LD1bd8umaG
P2O2BrSn4SRvJFG7gG6uajd6iyceMPtbcoD8NIFkaUYXWTr+F62+dDjTKk0fMU9Q
xb95P1CZu7v/kkBPXMpJ0WqQeRPVwqlqJjykSe24sRwhnD0nwp9MmS641aqogxFC
dwiwoW3Oyed7jwiuejRBDYWLWY6AzJuOKU5hDZbx+YDKjALhe9p40ZwIWRG9PjBx
GXJQh0gA6yKdkeXWOAfVWVHDmldnmHAytu+GSpLkRkDFKTmv4pzN3B6Ucq9tBL+n
3HF2DvgHqKC2/xyISRKFEftkVqu7B9vMjBa5MOe+AYDP6txY0kDFKX73M66/HqGg
hNapjZlT2qB7966GXcWCcVP++zjkSAVmKLoI0y/C6EfjC22aZ6B8b6A3Gh07EYMK
trNt0wRavVroMchtgtjIdIjZHnpxp9t41ZuqviVcw6GrxFSMu1hzD5zx9lJdfds6
QnQXPobR/57LvkrPaAHhbs27F5tBfa8We9f/o9VUi4I451eCX6WUZRonRyMrH21p
qrmvYWcV9y0zDH41ltxTjUJNFfoRXZvt72YLe01oeDl6FeMXntypDF7/Z/8bAX3e
d5Ba04pGNLudpWFBsNrG5h+Fisk4g9sZLDSYNJGLwla7hhla6E0oJvQs/f1Xp3FH
gmeP54t2npEqeL44NoCYnnrGVg9QgLL9GGpFZcZ7QHkiOV8Uy0FUESdfjYjmKJ/d
gvytQTxfwitJI1burC58z0B59OSRThKurgpXIcu2bpPJiTY7kYOUV2JDom05gWIM
695NfeSp2qKHuuUQCK7qrcULSz50RNRXVYBtH79j4dl7UAvX0y9IRmBB24YGPVnf
j+gzXeyrt/Smafd09OkyNLJW9GWXllP9IEJwBwijnpVjC6Nr3t3yzr4mOXrKSVLU
ODwRHYdBea5SJKFkHhw0ggQ6AmxvOhvOOOVweilq3bk56TIuzy6rgWkqb6keMWrg
4EJvyvgxVDkPD9FAlVDt/whZzq/VNn3IgTdCRZj4swyTgSdY8KUD3g31+PNNXzoy
MsEChnTZXVfGIJ6Odt1Alm4YPv0mvTPsqGKt1UUO9xpd08nxebElQ45b1kIDG3UM
89ZlKsCqUeiplcfUgyidH/1IaO1LcaR798WpsL7XpV6DibAkW1zszGvwAZ4SHPiF
Qf3B9dmiP5iImQDwp9Mb83oMrr+P2S8FPyk7ui3KGMV4TUOml1o67fXU0er+rJMZ
kMYISTCYJLCfiQRjDOsXY9D0c/UzaKxwyWfnJt+7hMvz+BlbJR7XFSc0SAyIa4ln
xweBi26OWe4MFn6D2v9Vq/KFv+bMmPAuDaUPUfbN5ItRLoOm5IkcfTY57eO2ZkeC
N8F1Y1shfM00klZR+B4EWDh5dsNX+epsZoJz0bFeed7BIA12PRaFeQexf+1rh8RC
eUr/+/0drKPpxj5iB7h09rF89SfptYvJpuXQ/J+mEszR/zTSssClQI7ob5zBq4Oc
7OL3d6krrEgNwzU0TJLxyMiutJKpJU9y+7OFwQDH0HWmaKMmHMkGITmeXd5DNmgo
+hWpIFANMYyVCKcP/2wysdBB4pvqidGqZM3HQR9TxD2A9baIoYE3EupDDhMJM3Im
qbIP7Z5vK3bndU3UjFSpf1K7OAVfvMJC/c9NC7CAFIs5EICZn3WOt7Nt/21qlg3Z
5XFCiaYxEhEg2s6XlUz9BHeYqqA7pUeZeAtIcTfXTngs39mWspXf4oJpN3f9cNXm
EDIKODicZL/+TZINaGym3vGpWGeyUkTHYKDh/T74Cz/PGJIO5kHqfJRNJPaKcOYg
UAGGW6ooiecZeP6dLfB8Uxo6TIkYeKgE9fPJYkfbN9oSD7/W/y9Dpy1eCcA98z1/
Jp1DSi92p/7lKJsOuBVmLXc8LSuaKmKUwP7C8eGKYBPSV9HlKCWrsc9nNrG9ivwR
GjgbFhSrDiKwXGeFngK+CWgCsllHZFDsAzLlV5JO8uNF5qEeMUelxlFQJjhnegnF
CyYPmrGIB3iadcmotwzOaqsma12wYISj05FYS65iHyHnL4se7ni9BAf6IMp31Faa
EKsWLIBIHOmzTCgxe+Q4hHcg5SMsJDI/5LB6YczFOe4JvWwthW1PwP3U0TY63QDp
5xrhHMYzGBkJnTc1UcteYtfHP6NZbVcLk2b/kCGMrft8ZkJalAL8qUEAiN1rpbrs
jIEYXjJipxsExoV8gjBTYMgLDbq/H2IvnFYXiTyGfy8Ej5+XeuJ53eIYZJP6ueah
KzCx8Eg9TA+azezeUuvH2CkR40HwmpysVyj59a8KbwhfuNCXqe68etuJd7V3BsDt
asSvXnF09ivxSPxl+dw2MpmDDWLS1F9gg8nWVLhA8CICLZ15xbwQjSiMH2KZyrru
ahhisbqn528eDAm0gfZFhldGDrFGFo8z8wRLQDpZLYWLDCOgHabe/dzKhTUsY6NU
CLOL72bulofQJmKhyg2LB1ybYg3vXpXF+8BcVF9K2RxDnNoj4S8edS4z6E+mUTQx
c0vMvtHpJzQAppLuXaDGDpIj1UxR7qVis7jcNhIEcBs0ilO0NzFBu7IBcFXcrog7
qF7ssoETEsLtVfxFyj+exFbKYbeE48OaE5zTxngnHF7H/fcz2py7f0Fm6+0sAzt+
nK0tM1e3k664maX85xHwa3fOOCR7sfOSpLQZgQnDra0V42721VRe1Y6ds8Z91hOw
SAeyQOdF6bmSmaGRnOG8SUjQvicx3XQ6n/4QF752xy3RLc7ecV1Q6sY7fyUKXNcW
6VT7rzJNKIdm2XlPGmdERs1T077ACUOLkz+D/PoealDN1KDzgtNdQmt5olYw5Zym
ZEtXrlQwGGucCO7vEJxwOvCgLF+EdgfXil6vTWE/Tf0=
`protect END_PROTECTED
