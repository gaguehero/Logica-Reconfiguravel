`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1oxBXE9Wp1EcahgYhgaVfY2JvA7J6oxIm5bVLuwzoYbOAwiNR2CDBKG4mNqiiFko
CxEBrFDdn5MY81b5oxvjW9elU+TIL0spfdSArGigye1883z81AvYpM+TkXcf920T
Rpx1EnQlZnpUDMnRe+51MsaMZwKgv/mSwa813oTqib0hzh+77V05B7f6d7RkiMil
RQ168Rt/a5qNdyM09o8yD+1HKWZboY1Khxm3dj9iZEJD2vWU9jhsNMXXsfmGbIdG
f2PfnIkaAd8vS8/oK5vjoSMmMGaXzrQnul+zQ1suo2hBdcrPV2Q8Z26lhCwKdKbB
F4BKYHFnG0GbqGw7PJF8XEYo+5j3NMwluZQObnel42oSlHJkv8IxMDCKiihYzowX
ByQ+NF5eUdTGOUvB6L05ccwuY+emfhJlD/pOhgE2ck3yB908qEOTaeegjTwrossv
AATNzbtF6GuNvXiokPBWCa1YitxRSppU5IJnz3UizjufdpGcUG8Rc6CVjqtBFq80
L6KChm71lLjQgMFy34SBAHI43sRyOZvJJjq8DEF2RU4orFGlyCTduM91QTwVGabL
9o3EzAi+HXPmDDTWjMgCc4WoBVqrQEo1vcS8mlIOGS/wRhXDE03ojRUCOytxKYPJ
J3iwdH98YwblyT1outgqNU6WbmsHo2hMZdDwL9ciNsWOZPj9SvjQeCjzKLzB9So9
vBvL6fvTGE2CYRMmr7gt9UxZzk+Q4XNjX7gXfD62PqQ3/FaurJhQtdOrffQL8A6+
1LB63t1RPIrEeWyqTH3gpXccjoGcMxPmBVzjdF4iXmZ/gjGH4DVl0aUa7kshj8ft
xbISXc+3eF1X1RyfjpTopeh5uky/Jgb7oH/bVl7rzUkcKp1HzYwYbWrB6GFYirGU
dlfhrx3ePmeYb6NWMk1jwdyUWPJxtfz6gYa4adM8IV0CMIUqhIczdhJqvgtq3p/k
3FP5IOvW4u+fJ3vLZuGhpdyToueb3EAaTR+6v6gqCuq37Y4rYdGcfvoEPxqPSAMf
EJD/s+tYcmoDJqi2nRA2/yESSVtHsAQ8q5s6pA84llCi7TJu0hypAphv84prEKxT
39jHLqNrPpShDa/PaCemQERGTMLc/a/SYUj2gjkZX5sRLOYNhAq5nuqXVKjSmuh9
jLRZS0s4iAgpnFFa9bS9SQi7KkwQwE1EHTXvPxWNDxqOBPkc51fIA5X1FEWYHRmX
rAEY/VO0JAwN2SbSLUbd5D64S+GXB+Tkz3THuQ95IVBNSOFS2FWisIP1ymQdaiuQ
6YNqUhwttRNQ2wDVFPbxM8BeN95HuK2ik6MEwigqgb6/vSETJYTarC8wNtcPZH9S
ZPkY3Lz39b92GNz8agimjJN7gYJYS8SrCpGzrQsGW67Lp0Dww0V8lqb/AQUUTfID
bGL/5ul8snBTLkUPYVwbGjK2E1FMrouvn1aciDwMCl2W44JZUCNZxNCXC/2JhX+n
QU8VEZFIHyVOjmFFBfYV9FDgMq/yOPTIZr5H7vMvnY0Wb9m2FdJdZ1/bmgrIogaN
SjBBfk3Nh6z9lz/LxembyLDQUnddPjzN3QTROPHCmentZ2aPR7UvpLY3bXxcHmMB
hjk0N3XNMbFoZU8tPEHHZJx3Ph9R8PNlgXx5Rc3RWxLGKuXiNuCxhFABEiMBZbnH
Fcw3RH1xX5dpgY4l/FlcqPseav5+VjLETwCtmd4D0tSwYwL5/qIzS1hNWma6J4Zy
0HSxIItQcynEsOCWFprx+LmWQds/JrE6hnPN3FOYNBMmzxvbqZHNNqIlnXD/G0nl
lYcHwgzCLBKnah9laRh5NRej6IvcbUdJJ3GsigJC0T3Q2G2XYHiDbQwuk+dBPz5P
1JCTRh65nbVwGZ3hLBYSrtsbx98DELYzUVZ+Uzhfsu6rdqJr1nVJHc7JYy5wJ2QB
NntZu/wnL0CLytzKXs6g4fxmAaLLhbbJqnFw/dysZCRRk+qmnRYJXVsjPrzw+rXE
cii+VCkk5iuwYa9rwCMyq+SwOBpv/8XPW/R/rZlM+e1BrjeSt2oRqx6ffUU5I/7W
HmozHLfAVhfuKXifZQf0B3pH6iNc2eJ6H27MuNWkvhygSL5iJzvpp7xxG3aaiGhS
b+KdDLK6kHXhblBeNmdFIdRQs8B6kDimIVgZ+uGejguFY4L3y1czJdh8uq1FSW7q
o8T4cVpXINjYYJuGv11662Qk/4JZpBh3qmUYfYI/+Om9f4JdcZenm3muxqf46x+A
CAzxKWgJeKyCSop65otGYZCEEbq11GKRORT6mzp4Gmkh7i/S1l+KU0NSW/fl91zm
ISetJ+tsfv7JS1w1/NXyNzmY6S7Dn4QL8a0/4r/9TehulWartegbyqu+F81i3rnU
jUYxQK9RKOhpxE9dNxPcNqUgZV/u2CLBJj1St/OgeZT7KeCaDcD4lj1sUa2QjYjm
hBF7Fq7w6Q+zwxy1rjQ9HIkLiVpP9ROZb+GxsKqoBEpeoDzRSEmRH5coU40jy9Xj
i0OvBBTfTjUZA0HY7qlBQXHLaCJaT2b8Ru8Hu83npIaxriuFvRQflTK8dZd0dIHi
zL1e2cn+y9F3Vy4sifUyXx9AKko41I0yutJMJpCm9czdMNkeDOfdWj6BDHV1plXE
ArXbZ+7SRYUP/lAEWJ7U9ENPueHn4wTTUFK8CUdXv5rOChyQwyMQ3BNVw6MzvTUy
EqtO5232HP+QkmavQljOy9XRze/ZlCdhoHKpYfLf1vRXnafcpiWCYXAvIVOSTgQe
AbyqsfPfVYgnklYmdVCiDPuZbvzGcWB5ovdpxWNXCeXZQzCTF1XTXSjwi3ZCfOgV
eK8oR/sDG4h2Gmp0l7JApNb8kDHedw+7iYy1z1iRWR+7NfGdNBovAD7rHWUDddVQ
VPik3Ypoa4FF2ov9iju7fGLTWpobeUz8ktGKckVgQ5509Bpv6TNcmYkupqVgL5Uv
U6K7AAJM6m9H+n3hUhVzTsjhviTVJ8JBwYzQK1FUz4Ba+tYhOSEkxyoCcEsDwPEP
xAVYoDI/1YMK3NY6jPmKEg55kOTSrK11z98gWY7IHdSv3JvbHYoDZMOhs6T1KGr/
nd50JCqHP8rgt0kCFRDUSnKtR/+PYhnwY8JPuQC6M48F8tiixAPjii5RVb4h+kHC
PeXE/LzabGY/y2GNw1Ej4kiotdTMbjOdRXghakWnHtjKDDWy18OaI9Ow2raeXATM
zruSNfEIkiCv+ivWm95h0zF1UfeLiLM1DFCK2KT3725o5BSDHPK6BkTLDgqTLeRb
HryLyNmsxkID1dp7lUv6MMKiI6uHqkJZKQPoCJZiMXlcs39unfBDNAzM5yTYshro
LxyOj6b75IClZ96vy1Bk2VSh7gFfpQYsJTTNlUZiWXFcRf49rgO6AqoAxzrG3OM3
taUJoNoLwD0VF/lRFLGRCjb2MAIhccJ/QhRUAI26jBOsU7mk0VckbiRgwyx+xavy
v6VL+EdWiOC5ORjgN+62q9ieX4PkcsSAToQEjHHaNlFTaI0GHx21IlnwEUun+9u9
SUN9pTVeOUIrSwU8hY/OgGrKsQJix2sQNpJ+b3r5sppu6w+gFJ75Bn5rCjg4H5KG
TOjnJorZTZMYHuYI5mcJwOFFCDQAxcJ+OcATWwT1CiL6rQ92g17Uvc2rJHpW8i56
j6fsvvHvC+u7oNHRAwYsD+UQoiGHa2iQuF6T2/x7ctdNzubtJnhQeLHbGdx0BLpO
rzNvCy7FBZTyCW1RN+68EmBPTpRuAxXiljLJzva+bOtNcfuwgolUB+jTCm8f2TNh
mQ1Jgka3TP+8z3/24GMCx/Rsn2tWYNVogvzTtxVXkYrogTxEI4OJcdLF5R2Xv91X
6usAfnpzAK8c5jv/I6rehgNmDIyw02fVeiC2FirBN2kbPTb6ZYYTPftDVe4xdPqT
xQsex4tnu+BVi5c8F4jF8Q2nEaV4RxxGa5hhoKRegxs3owB++kQBm9/kZQE11HL0
wqdGb5Ghct4hr04dEZwH9TgqCMvXD0uLfgz4N/mVXOH/p+lZ+QzVNnbkqDLPHjd9
OjShUIOIlglFK1XqCZh9B2xnU1KlnY6fAJRLNUrEEmiC9QHiZaI2IVzoPZgGjzA7
n7FazbcuKXePsV7JejLDDF855XCmA+qbsC6XeWj3GqSIgbbgt7CDQmAw6M/g9z3H
UIJDD3UK063/KnsPh59UIZ9FwyUY+tz0efgkUF/WPBUC+YxmdRNcsA+v1pCBcPvS
eBqx8WAgCJ0Y4hBzzWKOzclJ/ZNE8vDhQe5+XbDiHIUwi76Bkv5+OtyKiWUjJwhj
RqlBcm4mZoEn3QJTVJRsYcjEOA0iu3eA8ojvs50KdZ5D0qfU1IbkY6J9Pd4hNwuJ
bM4slKNLmAvbu+iiOGrQjpLZndFqCLqpDBekwOirnFm7kMfzgXdscOxBslIZwAYZ
CF65BiOTjo6h6moaZvObIMR8b+81PewSHo2DSbY8fQ56s1u4vJ3b//pcSoCvgELo
QK547GuwaZDnfQ5eE09rFH8wAzDaCXNmv4ww3h23p6DziDs8tlliuf2dumppkkTq
JhoXYnJ9B5s1S1/HoAZ850fmAoYJg08SbDm1O15RClsJtobKW9e9WePTZWVVZFSj
TGTmPA88qDUtnX/H7TVRAbol+/ra5pLzjYMYuAqWBu6mMxBut1+JSgOc4Uhzsqe3
kT4vxTLYAC3ITnZA0D7t+GcDQk4HUGgVb1fr1DMvV2ciEG6BXT45XIyhsM5tNQEu
OWZywXjAyl26Fa5cgXkbrrzl2ezecj1iBahppUUDBRIluT205Tyo0Kc9HFCIsDkg
e1gaLqGG+k1GhoF2SD80dZTGkhjLU0dQJ82do94asYXYp34FqobWc6CDtRsksrGB
fdavVY7Lvj0TApqFkmlcSTKn/8NGw3f//EDDs4iErDJvZRtelD+zwPovFSFDCik3
8RitEph1qcFEzMGr/x0o7JnWc0TqP3qru9G2I5uMk9BTxzFnzlb0gWSWwfZyZ3RO
i2aRa7N5HKyCZFeAhz9b+ZSkF06NkdD9/vQ0aU/McoBtzQ/tgVP/JW17GvrB2l82
bqfMNFJtMMYlDZNRjTfNF4OadR8aMqvAU0QSGytiqVPB3xSFOX4RvZawFNxfkbwy
Vcap/ooSUwnDpdJf3K5rIC603ziB/TI9LUx7t8cZZCwlJz3hhEtH0Xs9Inwbtbtp
fm0bth4VVrf/mMnYkA5lJr9tUiRHQa8WdWj/Np4q58u0r4va1nz/+xgoUy2nEeKz
t89KnAEoLfPW1Wv2UlzenGxgxPb+cqR+bwuLkAL8+RhLbfP0+cnbanodJwyunBnl
Gr18sKVF476bFEBDjXJv8gIwS6gmdY3B4Jzv4p219u/04fL09yqNErdDI/myqCTg
hg1nvhxVD3+OJ0Ox7R/gqfsnzQ/8ZLWPFQXOkWUkgYDyJrPAO4HGqQICieFaa78w
mA0sFIXLk7xYIXL8TskLZMZhClZvJi/Ie0DSGTekLCpXa2Qp4Zj0wvKsyWeE7iE0
Hp3agfwKiaeyLuwmcLSVpX09moDsQR4n1mNDLUZqRgXREOjnffoRC7aEQxH2PZUX
vMW9dNP9yg91FLQK/dvScGo95yInnxwDM4m4kK3RrmxJW45yCc5og2oCzNF/48bj
eWQPTHuaRWGxlDaFeobnrrgmQQadWBez3yrAw39MqXMi1VLYDXIEWvvGXbuXT/PE
J6e1F0koUWOgbQchrAf0sUj1lxLDvI4Jo/b7VkKR7JKI+GCAH7UqrIIK9HzA0eGP
ooM6075g+ttyArvXSGI2EK5eT8ctkbnSqsJW71ns+gLRhHFydx8iyuPp7aCVldFa
Z8svJL/yauJTlQVq5LGNU+qLI4XNUjqUx72C221RezMj3Qek/ge35Et4J1+7m+fP
hK0lkfNovdKAoGKzIzGhxKYEMYJVN+jg5lZiKHJEDpxlmhRWZEnJw+kezI/jOV4c
dyXjNUDbtqIoHyyUOVEm4mdiWJobwLAOszLFXJV4OFNUlY7YwVjJBu2uDnrVNxvT
PNPOI0JqezMP7p95+J13OdXYYJwRdFnNFZc7YaRESK9sLQ2gzi4zJ778KvsxT+tV
pJRPJcnegK9gkGrsx8Ube3gsDM9C2zihzkl0isiLmhTx3MPT4+1cq5EI4IDjBzMy
b62sz6ebX/YJVzDNet9+JF4b8EgiBILh0dw/lUpgHtAo/nsMV3Cz8hY4fkBm+mnX
Rsc6qsJnEn6zmqZfYy6mMmXiOLgdGq4nlvPYYR4aZzK/U12ahXpMVzLrskIm/vku
48iqV4+wTjEZSENEJbPmc3t0PRIVEZXcX9OnW3MfD8SjKcdjsE9TZHVTzaX4GNy6
igFCXJkh7tZTnm2E5wan8FP2uHHvlWuw1O3m9f9bjmz5oGoyP2mtADwzxteV1Cy2
t6lZO+lPfmrwjRsOTW5tCAz4oh1ogQLMFbA5Bo3THTVPsM9L/O+yspUFmTrOgvCM
mx/EaQf6Fk0wlsS99bYt8d+P75gxo59gJ/HvjxraSkn8KWslvy0iAk9cwLfZhDYl
PUS/gZMQH3/JLxp5HBnTBbPz/v+o4RbC5FAAfLsO4AfhTeVtTfgS9Hw5ab1k5LhQ
jPoCbGADooCJwU/oOUwif8UZE4b12CTgQPDzyQJzex1xOg0rVnxzbm795EkSeoKB
PIX5vT+KDO6l2myOtVBWl6WZSsjRfy3lydtqUVcBRZw=
`protect END_PROTECTED
