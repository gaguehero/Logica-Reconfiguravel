`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3W26HfY9UMC8G7Km3RALdSC5gkPMA9/3u4/K/xMJOZ/7UqRw/fR9ZMmL56YpYLb
w938ShLUJQhSQ1PhhUEuNWuMpZl3ZmZW+Feehpa+F+gh5iUwntHAL54bWJtZJNGw
IgLV79fsBssk1u2i1gtqbEw9EbNs+2+7H/RmhtR+vVdGmMWq3MhZvRVJZtZOKUjE
0aDU+946V5IyGbRZqQ1swIgCD4Ehp3ZjsWRyqSO2foTHW7WPnC2hiGiGULR+dfPE
031QNL6jDovP8eM4eudhi9fNrxDBdwf11rMWoRw5ntYCJrAkA8QLRbCySvN73SGC
Pb/dZDSFToBeoW6CYW9Cl85yi6vezHTaVhsUU+O56RuukYFaoA2m9Ee1HhmdpopS
5TYKzAUMxcYCOs2nGojVWesVyjlxKihNgP4Jwdt6+dnO6/UqUbeAHl11rcQmwIJ8
Z4591YkkFign5++XXrqhwYiggC2vJvnENHYO1OjpkVNJAG5l1QwVw3SfGX0au8D2
TSC3MP9yIH/3kIqyHrsnXMQ5gSr/J7iF4IL564JcMdS8dnL8lEVRfYCZx59icw0p
ArB33zJD1rZP7wobEnujqIF1e2dxzJrhQmTz1ENPcQTLX6vyH/mgy0RJexwIOPqN
/ok2lXVpWkewmw/SZS6TwPfCBuXiaCTiY0Jg3xkWQcglzW6LAMTHSpLp1+OkJ3uy
NqArzgjy/SlkEVWAvKmEGtXjr18R86ni+/I++Ss6xyRv1pv+KY7NB7hj0trgzsvB
6R3my1pl+vNGLu+FeLcjDYDBrv5yx6oY6YyNRX55apiHhXnYBoK5u/PCnxYGBdoM
7O7AyqCEUdv7Q+kLfhWnsGCoXOzgWVwIGcjGDMOxSrCJRx5FXDS6qlkBcQacavrL
nHU7Vrai+Ym1Hp0XjiuByVYwfTE1C3vWC+1hu2Haa9VCLBZGihu04RutSvjDqj4m
r88oT2XKqHh8yFrIDZRJKd0/n2n2oSLzxBXaAKMeCvCs7WisIxg6hPKbdWDxk5f8
BtZKLe7pp3Z2Wh1LA+0uYG+jUSh9IrrkPku+YwInUi/ndc1SZGIrk+m3XLGZp6Dk
NWgdrg96NbD9JSAu2BE6GzeQ+I86RqlfM0kd9jvpRulKDRm+0iiqCx7U2/5kGaIf
zGb/OgjguxlA4N9U2/F5rO2RpC49KrtGf+9sRCwoQcAwQhkw9a6dqKCzTvhrAYf4
DVw07Vv88bLPvaXihJLcaOvTNL8yVx89grJ9ZMSE13vtMJofLGDL5XnqO5p6HAAP
LnXUtjdPpi5qSO3+6YIGoYzZV5nDZH1FdO7Gh3TQqOWVnJ2sDHnwcqg8vloevzr3
bggIYvQSHZ5NfZqDv26PrzBKgPqwZ6RSOwfHg0tAhSnz8yn3hjV/RysaOgEAXpNO
YPo/+iKGlgVDmV6KSKNTndYt+OC1oTOnI+g1wUx1tnb/h8saSLEjzQFUO6hvs/Hd
nGfipc0htRXqIKTg8QuUHo1ZPt8E502CDIBD72xRfLXpsLSupCrfQuOMoiqLnHIb
hEp/UuxgiDYwIcK/WeVk5y6bcZyq+zRSEneLNClwM4pgdf8S/zHMfov4aXk2i/0S
pwdiMbIdum1Qw0y1c5wn2aG+bC8E8d9fhuonfdjAm+65wT4RVPFO37uzDMp6Ggks
9OGkKNhEs0YjMFEgxkBpHwyQ4FS39tL7vxygZ8WZHuPx/50yUmXBw3YGdvad+YfL
XS/izp7bfaLqUuHL81oYs5QXZ6IbcbbywpgqrbSH4vCEolro62B0kAyurFao2rY+
NN/n21goyqRXPaXl7b5UKIF3I1xadgz8e7NIiJwPHBh8P267wA+HSGrjoXu4kO0m
VsXyEahqLYQAi0apZmBwdczFei9G31Kg8q+mm5Ye9tbL9CdzuA9WAB7Nucq5XbjL
5usBvbpxGmdKJTypHkP1OQ+tXzOrHfjzI2umGtDGNc2EdH73TggKTPT8AM8UWceh
mgGJc5XkMeBHj0zyaEV4bD/kx2oXR8gkS7a4vtrFZxgU8uTg44MqDZ/3FNZzkTuY
`protect END_PROTECTED
