`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rU62Kv+WTsJ7q2fncQf0DSTmXTHluvNK/GO+6PzyZFJAeWbQ6isEd2CX1jTPhisX
Rm3uz5dXLhx0cTaE+xAe9YoM2kHQR5W8hnsUhFaNbWgYdemMDN97olUtlFDzk95s
2s72by/Tar0HxPGMwSidVCyjn0jn7Opa5Puv8rMv9Q+yjtf6yDTbTQMjFWFLkQOM
7hi3rs/4oLyEmjuTncD0PN7qzyIyk3DMMf+DR50z1bzVPBSeVsP2ZbGdVxR2PIEO
Ayu+ss/hEb5CTJob5/3fA/CyViyp31BurnbWP8bVEHLjYyc+sx14pQn77y5wIibF
miOvw6x64t2FthIAeiztBpvFYXlke5Zg662SmOPNlg0vbSLxBc29YKlhI0Z/WkkT
3hBrpmH+/i25gEx3nLIFsbUBooKLuMkvqFLOBkNmEzvzT1npmyN/6GV+bWRQKgNI
Sfp6d0kGOg8E9R/xIc7HuftdJDkBKNS0sHQ9MdaBk+7+nXnmQs3ssrjFi3oCeK85
GcOtPXiGhySscPY/vFn1TA8c+Mq3quIdYw0yBu5Juz6c8/8TD1+WdkhH9HTPRhGT
5dj4jpPcJqal0U/4eopAHyMMHzqRH1BWB5Pkp84c5srpHzj45fbi2FrXmt/Iprv3
s08alyZrym0FXSsAoa9/d6o1BJz/ORUV3uzge/BrO1OUyKKwdHszStkKAOFGPywI
eosjQckRmcBp+5bSEK3RX51sDAOmbeKhTFg2qNQyOnyE5/vcCDoVen+dDZUnBB5G
bxnlNt9BvaQsLqewaS+dgAQKRw7ZnSkoOmK6ptkxINZOUU+tFDt5d5TTsPCJ8dG5
bseLJvw14Bul1ExKjn5zVRf+yHUa9KOw/4eXEq1TwOGncEJUqxYHFIHpixEQ2cWU
qCke3IbxZbMCyNO5E4KpIktLS8l8qDw1Gf7d1+dSRdvwjlAltIODgvHHt5plhQtn
saV15MhSLkoH0HASEcBmgB8bED8rpBsB4qI6VMP5lBD6nLiFWps7aXZav2Fi3q4v
foK8EB1/Tvg/AcVDXqu2M3MQlDsF40wFmu9//9Ce6V2TK90LOk5hsjtwYZ4I29y2
lDfBjgsEiB1gf8UvMkE9vfddqR3wyu35fyvE+KhSs4apotZvXEu+e2UBsQuq96WC
afNA3eqGcLujKW3fkIRars+OWxcfbTiNxGw3TOazqMFtQV8xSanseIBykPhvycSq
MWeTtkpN77sEn0QVFX2KeEJQeAXreC+W2uo9VxF9Epqm+5mLfy66a0a4emv5FAs1
nLbg9xK+KqAg4EhCvNsbwAZRYO3NM+WxBTIvv6ZSc8gbT1tMdDCT3OJmcreDFWpe
7JywfxfDbdwDZit3dYMog+D4LozjHnZJcBCIzvpgdhGzvoJfriGyWG8dxOVhCAPw
oBT/r9h2UMSRGlq73OWUhdLq1BbSF0WwSM/dwwze0mvl9n+RRCc+6X6XEw8lWswg
UX05K2BMMPoEQmNl63KK/52ML1JfG6cwM0H57zw4d48+LaQ+yTQk9iyZlamgU/1N
b+my4OehLrI/YQIhlgfWAgXg8P3HGBT64U1FypdOpafGgcTXimu6gpScLcdlGher
47M6Z1IL5eRXYJ4T+08fH1WtehFkeHNTE3CcmGh9jOnbXaDsI1Q5bLK74GbZB2Oh
oHfYFklsdn7ue+hqcdx/zoaB5JzZIg5JUAxGpBPaLAaGOWZPU661s1s45g2QettM
gUxVovMdkTvg+FBbtw+54dcefMzTSxBgZQBm6pLfX7WE4AvMRfjzGwwnNqEGZsyx
J4jseSAoRPKpvvcSZRT3zQO9FBSMeHycARgx/gNyxDnqiZdpcHYU4ZkaP9xUvPsV
KJz0223cK+gGC7WLByVzp92EevHrg2Ov4Rfp95M0gg5x3i8PJ/fNcaJmKwg+O15q
QBCTCBjks0f+srBQ/UZW+1Hicl82aW3355aqdDL3UzsgN3ngFqzhxjTm1YGtuCTQ
+P9LmmoElgdcAhQfeb7/JUXH/VslkqZGyOR4p3/8FJTuFmETkl48WaK1jBA3W9Ry
`protect END_PROTECTED
