`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+1stDMsx77DNecUDBobBJgLsct2wdQHemS97SFjpaYXL/jnG8VpYvZjOXzCZR73
IoArGbxEc4NGTKFOXawNhpjix1fFXGChUQ5iEPFuQjuvgAsH/pZw9cn+7cKjz0eZ
DkVeGOPGuqM4xDwWnqeCMm5TQK0+bGRAfC6cgTg3Dmk7lTqWAOkcrzwPydB9kaCd
wHGuLz5oM7OXxoOLx3g9/NoQKD/pHuwGGfYKFzBwFww754Mv7zzTkuVVSHQ2VpCt
lsRAWPCO6Aa5xvZRaxUmuT1kiVpS6lMRA3He1KIJH1GBI+CCk+01j7dfJW+KYXBz
4KDq/jtFuLEuzLOEkGvPIrgfRTdBn/h5EpZ4f/drp/TucYfF3Qwdnpks1s0TNHtk
lBygSj9s1glQqx80gBiP9W5TZuzn0z1bZGID1SSpcX9Isyqcjwcz5xkAnQWqG/ED
RV5IYktQGklSkXvXrhKGjHJHBTVYI6t981WuTuw7GP9vpJ/E6N2u4lMnZojlRx8I
ICZ8U8/s+F0AohTtlwkLqwOOqOdmSgyfST8JECxsgktM9nkW91845FMYV+Et1lo3
9mEeOoVUhYdJBPAQTwWgptwgxQEsAhFWUsYPUShDAjEU8165yKjbcLa15h0FgAkW
j5n30Mnih82P9THghKu9Jkx/M2Vjf4aD8CaE35BAJBIWDyGBLkzkUaT8Gtid0hOs
T6xvV2zay3OCp7qmpXhY9fruh/pDdsMZFrSNHumLKDltOxgz+ZRBXhKfdBVrqMU6
Olu5BqLVokaY5U276vxusCTR/+jTxeZQROKmxFvVHnpleDI8cKIe463tv4cCGyiB
BAvcamJgkhxBU+ZPfMDn4epVuwoO7HBnSWxxh9xAksofBgd9W/As/XHHy7AFfZZ9
HcQ7qaWzyQdeqjdDCQzpb8/92b0V8IY3LkT3IsF7//4v5e4QQznVd1/TWyr65dk8
piR1Blf5BcvzgKLm8PCnAIzWonPoG7p4AZli8mMZkg5qqCogNeDHgbhU8Zpeqqz1
+VHPChHQC0uHOH8QXznp3sliBVXMEtnno92vllV9i2s8YWCmBi5q0sjh8LV4BKzD
bW1hDBc1F5VBy+dHOFd31SXkiPF8yYtSgrtjPk47HMGkWwGfzu/5jA9buFaVDG+z
3s38ilnVc6JlvFsFEx9AOW/JRZIhm5O94QqG99Ux6J0PlWkXDE8e55bseCZ1esXp
MpXUpMsC/vzrqKq0VXn2qEZk9t/3voWujYrZnyxLKLeeiyeSGm9OyR1Kpr8UKtBZ
m79QWMRIv157JwpliYP4TacFkERwbb+4Cow4UHmMLAdb0SYx71sEc0uwZSGjYLCo
q87Ka3R1mhgqH5GEP7EuoVSqRxSkl6EwjZAJApXh6xNkkk/0ELcAt6gR6hsY8ssu
x0p75/31HVqgUHidghLagKi/2WrpMszlUDPpVs9WaiAJOwqE8NjGjDT27LWUj8oo
fO4Fxz//sUNNCaqhK+woTvcpsbPEP1+yoxeKX1gaOpaAW/FjBSbzBagKdUrialwV
msK1gGRp5uGiSBasudyOu3InFo9RmH/ZLAeobT0DIfOVANKx4y5uq3L9M27P76+j
DEQTF4qL1KUrO9Cwn/xedt4xvJjdzmY+P4c/wGQW6NCb/McIbcf+Fx9q+u+nolXa
6+jXgd81gObcy45ysInzMTPqBKYLjqtPNtGJPgduVq00B4rGE9Qn2kjl0+ftYfmc
tcgHzRtXRWsQ2mR1aIczk3j+P9WBgqaJ50aChMcVT+UuEBZzmnod289go5+5wS5l
wS9KZ5n7MtK26VCvJPar6WinCvO6z9DSbgTQVhcntInmX2NOfj5ws8aXWYAGNlNy
CyUZAwoXUr68oWEpLGdvbKsfmxtq7umAgK2s0fNXvvcuWOI6b5TW/Mn5icl8vfZn
l9bcxZ0HHDRaqAc6wMjnZPT/9s06JAewGsq6ztZgmYfECLSG3Tun7HgH+ZfeTECS
f4aXtqY7+kpwSMLo05OMiQ==
`protect END_PROTECTED
