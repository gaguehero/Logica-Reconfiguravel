`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V926N1Cn4OAJ+yDZK8TBTbSPTEH5RzuwhSy75vYmAGxGECXbTQBfMjUhpQiIH1ih
xJbxSHCVl96dvnzQu71Z4KmSqYcSbhQNFFnaRCaGOBn9VUUJJwTNyUelf6E1g2Zl
AFpywGPgCj2iH6Eof0RIyJwFftmBdvAjOYPO7Gr3kcqLPVu/rc0TtYlpAeV1Y9pe
v4eg/J3FxbkrAchEZgJdoSckIVbDHZbjOMnCAeyr5omGrCmhMeD/uCaPmiM5G1yY
ne4ZVy3EIjVEVZD5wkEsGHoef4A+FjUSBau1KYchwgOAjoZO3CtvvmcA1jpfBPrX
rfaE2epT90AgNetpp15xxEtJvskfQG5nJVy9pC1D3nVRwa9XpLM4KYJgCV5FozAh
2l/frB4ApOUmJjH/c6J5J3kG9DuhJTVZzLBqzylQtWsooVgTYLPVIjSvX13CDpGQ
X1CqSpmhEPaAr0yLrQhQRslG9mOe2DxX8xbJpkpy/2QgrQA4vkMxXhSGWBuikqH+
88h/JjhYLtt+zCwO/xPbpjYs0c+m8s2o/LDTf+9vhBf01FtqwTD4+XGA6IZf3r0E
8ghHtrdvb5wcztVLlc/Sv4maMTxZ8zNszCOdXPKAFnYEqq/64Gn8vPbG4o+BCot0
s2ySAPwObRCymBD6uBhvggOIqrdRE70slXbqvPqa26Q2QPzPiujt+vtQ3V8WpapB
66HMHljrfrrrweMlvBeiTvZsy/DI3NSvvxz27BWMd8ZtMl0DLNcXsDG+WExJJoo2
Xp6iSH6VErlDUry9N6oXWialevU+g5ZbSL99wLnyWd2Alu5knz/L/KaXXsRqeLSY
UJ75MdjfMtqmJxqapYjyNf9hQ+0rIgMnqIGr0U2Uy8e/lWS/y82gpF3vtGMraCJq
MNScELkIG3wbcSaMOYfPf1d9l6lCG+9Njik1VrZS3JSzPK4v76Ck+02g+fhkKpoK
1cx8/vAKchL37HTGHcN91fU4Oxa9qLDEI8Rm+el4f5nmQUGnUYvjxOaRpDxhDxmf
yUMBxVz20y4BHCkSjzv6ubGnDiibPbDYCVNX6gXDVkWLXmNqJ0qp6aHeJ9rfCW7/
9G4kE1U735E4DTc0mzrcuKFUoTYSKCCecLogc/lrG85ev9Nt9aGuqtrSbm1gEXig
bfxJT+W9UwfV3uF4wJHGfO+KjFkDT+cv5HrGTiHC4KoEzzmmV3YzbMeJnpGW/UvY
8xPRzcrC97f9eKbaKgKp9/NRQDlp+nSk2fkL4EMKRohRQnZJv8fjQ/wBIkYVsfPJ
34Pgaqr3jBUIOwvDixpZ5/XUm9E+EjSXLlEJ4C3FqxOH44jPMTOWeqVDrbliQsqB
Lg7cJ+UgpP0SjwrknHJONTpDapAvUYC3rPtfS94a8V2L5Gf7a/nbOymPGf++Mjhh
vh5ft6Zb2g7dLwYUvzQ8CSTlpY6n8sjYSDmYSM5B6Ud0Plct1CdE17qn9KZum041
fMkYIItnxL0uYNN77hBxjWHdkclY+bxpTqC2UN0xlKnj4ZY/V1OFP4IdTOvu1XKU
NeR0YdmbwGAY3cDEhwYx6Fl+GOzFSZLKflFfPR9UmHY1gQcHn24DeRqkHjfBzN98
W+CJ+PUWlVx3JtmbMcocU2ocIcm/MViaT8kYqbacetG2kpIMQer6cnDL0hMTFGPn
KC7iYwT6UYcahVwmsZtCMZyl4nSdK8tHqD9ycAq4I6aFbpIQ8W8QlNZNCoAyjIwU
LCDSwSJKHROwXAtscK1sf+4SzqOvxyiRvta/mohc49VA8NgnC/9kAX+ZAuGXDR0N
4/0BWmACSuUY8iz/hEm7bTuTGqkibWp98r+ZXUfG2lAe6KS/0Sj/oUYCwXBIf8L9
lK0/gyqzI7wF9IJi+9WbORL0Z7mNDWGPYPad1hGffGnBmMaf2LAaXotOUF+fDGIf
4/L2veYrwAHjRfDnKEhHvkrpW2ppDWXRhZeaqRqCDdT/pR5RaBct1NbScD2dkGLU
0a8wGXIIxJMNtG0jNk3V7lYEzZ+CnvpcCgbyz9oPhe109/fk9Qwn+MgO/G0XchS1
8iWhl+AGFaga3FqwkMw9LjluU36OOSypGfgp7pV9TedcaBZAzz0rPWCUfk9h/zvw
8sAoQPYX0nqH7GaRjs8Bal0WXfhzeU8RjUXhNjpf7afsmRufe/I61IF9DOqVeyJz
E0gU/P7+uKz0eq8bs1k8KjknSRus6HlvRc5c8djnQUO08xQiJvx9M/Yngi9vERbx
tR8IGtiY12yl2qrmDvneZg==
`protect END_PROTECTED
