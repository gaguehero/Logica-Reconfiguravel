`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMhzUiyfOBX3KVx9YKdYHzON8TiPNz5VUd8mHFTzc1RjZHVE0+iixqy54Pwgm+IJ
eviFatRXzT0DGL5T0zepCnXRxkeYsZm3FmWX79DeLXkSfe2zGhYBwLEWwn0SeMl0
/FN3dwjpV1Re6f35z3HnHcYScCoelO5/omnKHwR2d7vOoLQiXAVEl2N278RiXaTb
BM5dmuIVhpUzcsJv4gM4M6MRLZaH146JUIcsSOU4SXKZhaW03WNL5n6910SnGLhi
K63novEvwcVfSSTQh9y7FBgsSAtPVWEVRqKFcxg6u/6l8B2cpgSFkJpUv+bVLgnX
PHbcd8O2/iEiUBiua1TiT8xhQSHOZWFho3b68tVLRu9lL2xXfYLhXSkPeXlkFInC
kX39W6ODMukJyGwnDhIYbeFd9pYichRd072Wr+ci6/SeehllKvUk36c4JGY2R33A
rzv6VQBYVtXB77SHA1wRbzT8O/GYoqVc8F2pts2FwbtdHm0ePeSFp5EoUIdJ556p
agfeLSoKee2XrqIUfkdzJ2BPeMgmWNpJ2I9gAW01TPBRksrTK7TsDQyovVgSviv2
a89gj0LD6zY7olldk0Hcr7xnyneSgKy/yYy5g+QQXQPqs35OqJHiOWfrQ6tRK4xj
ejpvAAqAcVO5mrAgzbXWXQ==
`protect END_PROTECTED
