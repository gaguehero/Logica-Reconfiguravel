`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33rQ0XeDk8AqRiiYOw4V4SUuH7mCWLtYqXPV6IbPG9VoRp8ODAXMwm+DomkP3s56
yKH96BNcSn7ulh29s+gRASlcNBF/tGL07mZ2XUwxZULVvFuPVaDZPcndk/XxdMdt
L/2Mlne0xueHc9uY9PSPOiFXcCWYtMoA6kTpxtdoLTlYGID/IEtRLF2hS/0xbBDn
y+Am5XnIjrpATBt77mGNPABu9GU7Z5g9kVjeVUSwxpA0vawtMTqSlLszoy6OLkMz
8wPCLUUtZiLYACXtSB3KJrAhN+oLnVaJu4p7EBsCLqB2wco02HO//e8nb8EnENrC
/QEt/s+Dt7JPz091bF0DUBAzFyszkdpkwXqCCLnXZDd9/fkVYcwM1mIwOTe3GUBA
D0PwP61qXzvb5vBEvblvx6Tnz2ac/Y3f3JxcpzrlXoH3YbWpp5RvPWqxTVLiQDCu
cclBex6IzQVdB4Yk+6+GQiqeVFQ/g0KWZZlQFKb4ach9/0lg8UyL10CqSpBI8Iu3
MsuufeU7TFekyFPs3aJpyJcLDmdd4OUw8ZpimGq5PxSS1Ypy0jCxT15EZDJMv/SY
5vtTWY0ogAMPCzd85x5CogvaHiguhP6Bsb/gQaFY2wXISFerFAAqZ2+4wtRhKxP7
akkwqvoA9h2Sl5EOwqIY+OHu2yOVaBKf3hFBTz1r6/AodYN9fNNoYPUJysAqbSAl
5VfefjHp4T7J4/z3qgVNlkehSFuFu9215VA7NpxQnjB3Dlp0ssRLEfZqI4l5EMZ/
PaeoMB8xqUUnOrrTFok5UZE1ZYRfE9tWCrx6TTVm/Uz+21k7LQEAG1I0JMWH/2Z/
G5EdiiuiDDK7OtiAahni6ag9jXdQCbRpZVRHk6CclQji65P4YmPFZMjGZ36ejNCI
wdqNveIGR4MNavFsLPisvhS0auXdE9H26eqstMCAogCgN20rlNUMckKxgvVLkbHX
Bpr+1BK1XsLOjfsCOaFW0so5techTmQe+3ezXNM3QTuwpf3B9riO1yHtJtzskYfU
ILjiitpjFuxtYmEdR6BsKFJ4hQ3j+3fiOUyxuqngm1RACbo6nvgEbYYU+SlQSt7J
36yIiiuNrgLq+v2FaqGLyM5BEcc1VdwB9pRFkCqQXRKUwJH1ahNP7lkSj8j71jLq
ACqI4b13OBNN354gDRk9sJRkhuVCo0I66+AOlyxNo8nO1Rj0my5aZ36SqsSONR4T
hv7+Y82948ToUbK/6MBEXH9mkOAoLlhTn18/wQQK6f3zGAGYJZFa6NQyAJgQyRHb
Oz0DRF+4ougCJstRBQpK0M1mT6qkuytXlF7hCJr/fDVreqb74OeGTlK4YHht7aTr
UkhJ0omTvRBpF3ys0rITQjgOb1R1QCqfcWR/y0e0ea5cg+wD8jFqtD3DbWZ8686R
Q7bGum9fetitRBQuGCi1Yogua+PvhQ0TAEZk3PADngDAX0P3QVpTHLVwRlp50IFE
uebUKEQnmDuhp72rac0R3V1GFbwBAVC0aX03P3b8jSvCeScb5GVNnDyTrE88S1p8
oq2EaY+txgNlR9Ke9XGC9a0WbF6/gzDUWovy+btO451G8QLkKJCGIj3W1K5WRmlh
SNzx0O6EoNaetTYr1gPEfAr1AmCjK4TNcp7yDQ0ATBzbml2R8KBc+KBmBYBL97xz
yrYaiLID/aCRM0aXSBUJwV5+Tnqf1EpeUkKzKiJrq9H9qW0a5vNVuVndgwTeM72j
uIx5AlvUnox8YTkm2+cOkIcANAzNug1qUQhTe2wbnhBsC63nQ7wYcmA+isu4ClDH
QePCkOiqWXUmQ0QANaPK9FKtI9VJN/Hg4+BAzhsJa6I4XSDPmDBxOjTmb2w5b6V5
clAdoGaP45BsJzYcAMwL9h5dYUXizEL5VwYOQDgfJyCFKte0xHcKo4KyLTZ/ygZO
XNroRizhsrjehSDVmLbclC2KweA4heSUnvyoWHBd0cl/7Tqg6FkctGckJZ7SjnDn
V7csFV728T8UTs9DsEObgw==
`protect END_PROTECTED
