`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5BPwqeLHulihuIBr/G8/GSWFBwM/SfbUVl8HRaSOooDemcSJ0SKT4YDbtxEVXzq
VgDtbnycPWgAujF31w9iFRo5eJ14DDroB95abKSAuRzpKstidyrxfHBrCENR4PNS
8+ywkCuSXpIKRYrT2HX2a2c9f3nBXv9CxEuO1xumrG+JYvdt7XTGYXDRdYqISqHg
a/deJFhc0I4gLHc/EnzOt+EJG36tQNip+N0gVL2BqaADGvyubgc7GmfpdErD3X5G
SdWiOh5x/R8BH9xltiE9kk7R3TWuOH68BPpxQhHCDXSnFaIMMw3fRdtBgIgU7fgH
80eQ6RxGKo76SzXn5P6k3k18Cxq8bUo3pDD3ucPttcnePW+KY+Vc7QzPQuU+PjCf
/KmE7LfLUEaJT8XbfuXtqn7wAOkQq9JqI+WTEdcSljcP8GFT8JeSg62AO67cJwrx
gsOdAIWwUg1uuzJjuudP+/15ymdd0M2IrBygw+x1Q2nhXqWnP0rV0j7aBAWpf+II
2Jbk1hpelarNyR7J9RO5DmvMqY+bGcNPYkd/XiQTtme+rOYINsAeMwlymlzc2br7
mWJquy+R62CIU+ZQSQzjRG/RwzSuv+FpA/C3VN6XDb2RxFjJuGrm1eSd3O0mfABm
Xl+gZXpgnoEzyB7XzN2nsVif9HMqFmcGxR/itIwCKxGfmWT8Okr2R8jros5h93sy
mBY6vnPcpK/XSFTfDcUqV68+MI6UZOPG62/sa97SPBsRvpW/qGgU4iAYEDF8wMJo
PWJAZeEZGmIDDF58xEpUbokN+YHUzauxIfFmPjCAGcqgCQ0xgdVPINmDD+C+dUrB
rM0r4ZmK4eC0wkIIXDOe+L4dlCUqaGih5Dag6+Qr0g1bZpgG228SBe+15Te/mQu8
/lyBFMv70uHkfzovVtwN4cITj82NmJIFz8dx/AgQSsmonlWzccFchRzI9+8cxcyP
YS7kDrtNUYNAhvXGnCQZCwKY3CEzYO8mLzYSm0zJU9dlO2l9D8z9RpYD2RLK27e5
mDNRUGiui/pYdkvg5FJZNljZZ9ceD41nzeW5ot6Mk9eqyZiaRKRL4OilgzAMAQGI
kvGzH1mHs3X6pLP+Oj2D0WbxCrYXBrLv6E+CFhUPgk4ndlrCRJW3KchL6PTwlnzs
Rpj/a+/RdIZJprtxxk3ttSyj6ABLDY22T4QPHBMf9Oh74yLG062G1U9kio7rCNQ1
ucmzKmH4rHBOqAVLwcMKjzBo+n+Li6iAGzu4lfD2/LrZtuIRZ6dP5fYJpycu0vnz
n1Vn/QRNpoSXUDYDV6N/XhkupVDkU8avaVyNGbK4JoIBqtNehLkVpS23iJzPrG48
bvn5+daE99cCa0NayNuy7PZjDrszTIWaOsmUq4d50EivSVtp18BGRmP929Wh57Du
7jDDc0PZOzrl+PIefmaZM2a3rilEx/yg8LQAUIvbleAdCzL8rHCDMjLUQM5aqlw8
J0XHH9zs/5ovw1PDxnpsBqtwVlds6j0R0D3OMSNmHRKbAyXP8ebYPl3ofVUrQCXe
vdOOrBPThM89ec8h0JXTzAF4tFZPlvXaYB05VUSXA2VpSgK9WHGX46Vl2de81LuK
Mi89A9M8gHqLtG1LimXPfsNJOz/oE9aP02mds5YAyhNS6TKTmeRv9aK2olsfMogz
VclUSseGjov4UlQShgWsm1tLEGFbmQx892JTXKJpxqqjqGzdSGZx0tJKeG7awhDL
wAF4VniNtGZmRUrcvHWlLUKmzQQV8xRCFioWWmLdIw75wytL75rgLVgqqnGUb0iY
jwWk2Fl1+AgiIKixYSUrKW1EN3Uco/RNfc6rV3GbjjgFo0BeSq4LN5ZeUNOZ9HQB
uPPKSa9EiGLr+QVYOAKPkB3pGotDluL4xBGzcLX9CzZqrBgsWreaGoE/cp/h4Qrb
8WlvcirGeoxsbp2uC+HuJzsssHkosEfwiSTL+CGrxuQrLhd2ygZ/NipzMbMRCQcy
n29wIRU7DQTcpbFS5wyVjw==
`protect END_PROTECTED
