`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCXi1KJIbHimtEbqpMdxSMPBkYYXZYCjw7NS7S2W/FGflIZj2iitqVJSODLXsoaR
Vr7yG+YZ+75yqkkQih9dRSLXAhaOiCTHEjleCSKd4KRpRL16Heknt2z51LQOscy/
fFmfG6gwWBTLQ4h++5xyVD6JjQyvQ4tJQ4FkauZ4Uqi45XU6fqeNvxC2PSBpSlvc
JPEvZOzDCp/Gviu4hG2b5mwq22tFjcuNZgDwla8xQAFCthXdQZMIv4yhTBPQq6jL
hAyCMj0hjgWf8HKqwUdzT1jSswdVBS0f9eQCniXVAIURRCQBldeN6exSoXPyUqn7
hJAZG4jb0gBZlry6nNlpWU2ExOltBqEB2SWrX3TZz6Fcc3+/krxwB9V9NnbpPvaN
o1TGuK6Q3y9WgvD6fqZe2RSiT4CmiQOYFNa061UDO/ss4JBuTbjpYUdaFpOhBsxY
qrlUw9PkiFeVzoea3o4ok0SIJr7gU1qrC0uTOJsvD7r4ogfhudfgNuFDEKfHNX95
q6c1TRmMtSnExkoumBYuEM7CWujmncqQy4Oppdf29AWNpd7Ldqbi1atIB5Q07z/S
fXb42NGQNA+NtRSq6C4IfCElvzRH47GlMLN4oadxeyudm8u4lb7oVG3Pp8uApsNq
uzzOtgP9hazXXdr3Z94WgZWhLSRtIv6XWp3PWNAFWJT7rV2rg0jlffhKLtQtQn2Z
quHo2/lcjk55jZoQI2UtnI467ddNaQp1kZEq7uGCLOYw/EuRfwSMPcjp6TyqlZRJ
rwg5bWMU1i5cEkNQEykbxFtUIr4i8ZOLKP6juPpLoUai85VdKC/9tREzf0MRwS9C
09Ql7RpIggewbZNGEA7rIk6ar9vxKbXcLSY9PhGAtFPL2AqlxOIe220o0CUmPm+2
nFklPUYrLMwOXYU/V6Qv/G7oK+hOOAgP56blxCrDixk5xjTo833TyGj0e848bjy9
3Huvwqi4uJBikCUFx7Bnz6atpqIrs6/qj3ZoOPnXKAslQLnGEr2KD5m07QKJPsB3
UvgbezzEtG8RnDMmhjYCkf9ZaTZngqYABb+B+oQHv+vp32AIgCQLNBLRqq3si9Vc
e5YQQ42MAAjr8pmn1hw7no8pAb5HIA0112TUU6UDQPl8Qp3HSqNhCzTtb6noqVpn
SnBP29dew2+sXuKpKeiI/ch7wGhfrBptXuFUonlDuiv2j1Y51nvWGfnwImaGUU/6
QZX7qcmT4lfJO89hLY381kPEfUsH4CXIF14Jb+28HEXbQj166FjIlNOMx8WQ6x/J
xlqRUQZqPDxTDBWooTimVm/xeFTvNgSUZG/robSf3el3+tXbAmhG/4WQRbW8DqMf
PCI0iwHmWo5BHwAoH0amM8HCTQM0pa1lTvHdItzfhxzBr4KulDhDEVHctFGZyWBb
nP+FV0kDygBkNXUaBGIUmLYhtYLEPqFXtZ/RcVnHLl2sOJ1aQMVZKE1woDjoP5H5
Z+Fr04++b30UGVSZym+eEXpoV83IPmk9p5w/+Qr9vZ5E6mclX9KHHDVVMmPsiVQj
+FeoIgPS6nuB//15J4Ehru7xXVTECwxBsDKdDkn0jD0wMdEfCjkexpCPA+ILqWgn
O1g8ddIp1eBN3X8iaOXFrHAT1kwOMN83GxSK+PpJyM9rDxIsLS9PCFQisUdDdxNM
YOps0+pIww+yNjE6m7pcnJQFlBrSsfMR6+EioshsWNZOlQANWL+4SnaZxtxRvZTc
ujRo89/lZNHNk0U6SYAuKY+HETMK2KJecDrlMY/YXa5E5U+gpzGeCR3YskXsxcnj
kDEIrPVRhvrVmEAsW87B1PwibLJubP1tXuBjwempGg2t2/vaWCqHmUoIy1khajF6
+SdQdXLJtjdQf/+Jtt/A54qkUoy0WpWT+8YcdQQJg8o4tiwVPV1ikb65V1d4ZaCK
pXhWQBKVUP0iVZi2slzyzHgSGMf6fZFBVs48hkqym4//kddZai+3gV6VYtPunBR6
PmQDQxHp0JPs4UZWf7bfridlInaeb+FwD4e3QCHmzBtzVs8SUzRXfFgpJqbkE3gD
4jgVtVuRsD5EDekifsNP/gzNQ9WPs6aoAtlJRQk5vjfBsx3EqlcK2ldnh8uxuhNJ
IUVesXkva0yoiOjruQQGTfEPc41H7++6L34j7A0ZCvQH3CyB2p8C0YAHBcZv7GQd
aSC4+dyhPTv4HvgtFSqPS/QrUcjKpA7aWjGdidSsUrUQie8sJg9SlKMvW71IH3Xp
Mfhwg5bAlgD98XL3PJQoMw==
`protect END_PROTECTED
