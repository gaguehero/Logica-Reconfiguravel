library verilog;
use verilog.vl_types.all;
entity my_and_vlg_check_tst is
    port(
        O               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end my_and_vlg_check_tst;
