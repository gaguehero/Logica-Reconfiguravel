`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qt59TuPMdkm+eVB/bIPqIyfhND+BqLt15wopbCUESBdEzGDVsATZLvCqA+c6aSTA
EuSGF20BcgFFcO9pj0k8wflvDUzPkL9i8DViF8Ka8Acr6qsLy8rc0ujV35oC1BW5
mlkku8vPkuskypuvXCjFsKgrW73PNrF39B/Fw0hYiDAAY9dgzRoDf0HZWVnXOAJw
4pD3AO5p4sHvUeHvNpFmClP6Ekp5ihDpr9W5JuUgl6OXoUj1wTPBHbFwG7W26M9c
SwU6ruk/20WFtQCP1ZZHkF38BqNkL0iTfmBHjeBIatp7zhCb4DOTAGG/cIjW1vRK
QN42tg9ktiKtAGl5fgXa8Ea5G/R3MbTIVE8YhkqW0wQMf2pTnSM4eTJmKPJP89xV
knjXD+4uZNxYIGwn5jhRx87bUYgY/DynMpzsiiwYy6F98pnaL+4WG5sEKMOoHbkK
tDXhOkLcWVD4dXDN1c5ESVzmh/3ZblngaSFg9my8szmmo3c1vCIkzQ79X7PWbGi7
oRayvnR73BLgpGWVEWm7YM/sx3EOBUV2LqQu5d+Fk5fCg2tdWnjoaG0aAaVP9DJJ
3Ct0msWetQd3+cIgVhJJznZI0EOTIdV9c7+k+YJN9es+CR8r+ltEjrtwU3kYh/ZS
u3ptk6QfEaCVaf5t6KWncjXmORl1h3ePFZNPAjwejdkdS2VQY80GW36R/KxYzA8V
`protect END_PROTECTED
