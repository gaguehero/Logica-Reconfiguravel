`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+EYA9P8rIKKI/6Q7d9GD+30Yjw7r7nHJe7LZ0wT4F28d8qU9+GqWh/axMbM56Ko
ow5T+lmzYXASGiSmpxo1C3svhYXCqKoRQ5EUZM4qdyfY/YGy3O9lyeAoEZ7LTHcx
nerLj3aJTkDHjTDTNk8DH9ViuVKJ5YvA6M9aOehfA4X4VUBA5y/cFvdT2RiOfiIK
2Yv9hj8amUVXquvYgU7poLoKtxaXPMUux76XTOvUNcvecijsXjTUOxw6R8hKGVrr
dRy66Tdm8BfTUTy92+nuLSACpJh3wK/Cgcfje5Bwjj4BeZW89n3rl1YS4Wh6ATih
lwJeIAZESiHbfchXxar3kCF2N8bmpbR7aStJeF+z5yqW4znOypdh7MO4PPZOHN39
DXEpV3n+IvSUxbvS9d3mdGQP3rHwkOizIKtjDiXdTVURmCM5Gf9imLr0zCMYx40q
4yQjsUal0nw8bweo0RUjt8ib9Fd1OGmmWp6+adrxdFpzjcNYaa7u5CTkLnEehjJA
nFeQZDpK6IXC1TAc49MFxn+TPPtQZQtSyvUlU01G1bBK1z4cqVfdxNsWjYsTa4GI
ipoEMelPK4vwWqefNTiUT8EjOunHwGcxI/+HqH5FZzm36JAmGtl4/Yq/Jq1wAXN1
hG8AKtEo/KGKUXjjwE2YQ70/yz/yxuC4oFn1M6GHrS/bjTHo7L6pb77dEnC5LizX
5VLx8BeiKQY2foaw0rJz6dR7CyPX24V7A/2M8odwR6iaKZcZqgYhM4L96nRfM/GT
QZA8ZGTW83heMqVb1Oxhh21M+Jp+kFSDBe5gMPTxerAdnPBfYSSpMYCMd5kXH4Wr
fYqOyTXbIA8+uFr52uEJn+W276Q4E5qDOC/Tr4892WEoPEevScSKc2DTBnRxtYXH
cTP1OhDlFPNsPIpjnC5d+QGJ3tF07JBX9FQO4moSdUXGdObIsAAOzMWTiTwOtb51
7bvY1xu17Ir1/2FmxOBV5P7OOD/yFpqvjRZXVJsAwE2qqXhhBeOXIt9OWkS2l5FG
iIDletG/+rIKgjuLRMvaOSWn3NkyteiuI8jefuMGwhFNxtNCR5a1kDNrXnq1r9N/
Nm/yZ7HT2HDq06ccsDVx1j90JgaKVF1rbxjlgCwSnXkQQ/lR67GrZrVUc41Qvj9Y
yWai619Jc6oBzMVPyWoPMeuJ5Z5AAhTKHOO+ff39WQlld0U8LUR9wAVLlqDxWIli
JOsFllqT9zeM30adJKaJH+7evNNNBHaptQABR7i7m8q34y5NmdS4WlURrk1lL6ND
baY3jcAcpbKDg2nLhwM/AGdR6KKOGI8EP2fHnKzPEFTnlV1GIhzqVKh1YCQQBBcC
VvKgk30zlijbtTmvup1LgafiM2giuIWsQRIF6NPWL8gFqvDtHwLXGaq6OA9+uozD
XwhLorWFd835/4FSR9/PwUdq4I0uLA1bp4JRcsZSarSxctkKwru80WzxztYwtudA
/eDwAXzsmi8efxAY7nVYxRuAXGoLYuQdK289uFVZSOH4jwNa47XeN0qd0EN4c8eh
f82cO/UTnG7AIqiAbYi6aioz8lGUfIMcwon2HmOJegdF0ZnIVAYNgbucIbDwkO6L
fdvd5Uc9bD8FLG5sq3gO40aVXY41yfWFKUl+ofu/q/gsS9rft5XEkZv+LIOUgwhO
VK4HezlI7GlFEAEagecIPJl7PMR6Yv8qXBuSe8+z/r9du+/YYczBndelQyT8RIcQ
PRpELQ/BtbpTJe1AaK4XJOif34BfIyJ9IpR9nk9MRQnm6+zTWGGkmyojZfTOfQl3
ALMPi0H4kdyIQul3Iu4hkBp0aGwy5SZVkfFaR2GxdMgNU+OatYwWkarVDzXYNlRd
Ez9u+RC53YudVMZrRaK78k5dYizfltXUF9JtIKiV2LgfzeXPBp3/CU+OZy7qV3mu
gVump8vdbVCnQ9YFIg+0KVkRHNBQNXOfqRf+C1bdkU0oC2TSN2jNr+EFHRhAA9pY
c6l71x0pVCOwMBvnWyXD3E42VjIZGi35KeCMi8zAXuR7of4JbfQ/CCxaI7i7EePv
`protect END_PROTECTED
