`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZhZ6uAcoinYSSYOz/lgVn+5J9TPDukasMQ8TPgywpZ4ILwPx0nue9ZSe7w3Tlr/
2nmm3RehhnTa960JfP4RE/W1hePFaWyb7uq4rYtbuqQv1DMIfpRPAamtwtPAxLkx
+JJKIJ2/pnfRZ1z3ndjkg8TRpOICBr9r4hNXhoehyEfg6XrbBErwRTVWgkDXZ1Iw
5b9amfk7kkJrJmJTDg5We7TEtBcKHg+mLUPc9ieTWqhZ2nQOkhFyYckNnRdpIVDr
k2/tWyDa+c/ORgeQjukWXAns+AK5VGnr01280nLEPWiQBGvIMy8NeFmFc4QnLG/s
LXe+6eeame19EdhBuLPS6dA3tpIuqC50SsDe9gqPQYc3UFJWzuxmA4RDlb+pRQsx
b8efVo4vD6fTAUtRXslfTWiQz8sdh+1OcsapErV0e8tBqzYQXmkzJTmoZSMsXNwE
sGXWvhhXttMRcBNEJkbj8UjjoRGHfsoUDBtAMemsWalNPTg0ha5OWt0jMUzv/T+j
0tR9LHJxoiVKQhaP0BMD5D0nBCaHSldlSGUSb8NTLB0hd1BfvQfO7JsfVnIPI9Y/
3gU0WlIAb10yMmlpzFESsZlZiJUKe4C+gMZVnMSD7lMDphOrEL1z8ljFA9RNUp6w
sWZ41UMpKZ7aqs3hJpGx7g==
`protect END_PROTECTED
