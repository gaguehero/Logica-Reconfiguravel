`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W75+mhWm9x2L5USWMb2VW8Vr/VtRFVPbcSlDNNlH2LZo94NR03TTMGAe7i4Rki2S
upPa4ScMgxaDDiONB772KELWnDWdDXlh8dP79zz/3lT/mtn5WbMN9Tp+QzrU0D5M
ZNT9X7vtqgTAIUmpisaefDOx4LodNm54lRSIljEr3T7uBO5tCg4f1SRLBXOsVxJx
2Gwop1wYqRjknMYdddhP0tGRRlixE9tBdTivhxgGdYO+pNUfiOmMPdOf8WEJC3l5
ddiQpnnqzmD5ACpGGuchjgBhfjLBPpfCAErKQSzKXR4cOMeOFaU0go3JeUqPKagP
FaEYx8VDVpPJnDY0T+kl0JpbqxvLVvrYU0u3Yo4uyNhWBq4FZWDoB5TXVO93NaAw
XoshENEgVXQh6X553SrGHSol4z+uwV7x5wBTsiPR7IUmHpLwxfCagosDjE3G495Q
lzXNYqXiwxRscxuFJwcRvoF6SQaI9KzDR6OW//fE8gfk5OkO/E/UbVHK2uM/4srI
XsrNRffvyvjtdHwebBUEGd3LzDXHDHxhcTAHNIKln9LU2uN4i4xXx3U9Ad9ahRB5
zIed25Pd6MboXjSYlxKWP7m7/VB/D7emRxTJvwhlJgCSsZS5RXthvl5mg7FN6bZo
2/Ph0P1nZ5Fbkff8jQe9JjlHSjete5Sxy6ZFyiHMhdBXGpAKIf+E46w156FGV7mf
`protect END_PROTECTED
