`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6CCSBmNFP8kyT5Oa1zxtI5tyOvYfShlrsKR6wP7uy+SRBSBIn2C0VXk1ymYTkhtA
QzU/SR1Vpfr/fFGgSmLMHQDADKEn9DiEgVjAibI65e0phWRD/fgDyRw5t42xeDnr
Ss/czTlLsr1DG2+aN6/ZLfi8YsUiOR9ZVLD9LbstudfzcRPfSFWidJ8t1V3phTBd
bfMd16sxPsIEJv7PJuwI9S3se7+oKC0G6ILpuXPpv4bpkGHdn3LFgiGx/pxCRkV1
VB4Q2GwvMXknZPlvTYUaAIbGkSzyw/Oy0XRekhV8FwoJLB6YeJAUlB3KBPvEq1TK
v8Uh2Zb92/zibfFPB7OXIfI2VgFb0BRl6NGqiAxWh9XBQJ5ZP2aT9RX5N2jOeyfD
xNJZHiSY+cOpmBqUtUiqTRwWiEZPUQgDa5F0FdpCk+1yFGZ25oksToOPEFXMsiy3
CcUaK725RMDr3vSNwv1LcLmouzcdBxMZiqJdWVtWWcVdsBYRCVtCYFKee3ef8qbH
ai7WGH1osNrnq3PXWeT5Iyh6fGdGPdez56CcWFjtjqdv5TfEM3GQ8M3CHg6b6XIx
LHRd3qV0VE3e2+pu/hz+KLbFLFCKb0hzn6xZXV2YPfVsXnq9tslP+xuRIs5H12uc
wjrkW2d82rnKqk3KhBlpOszzTwQuWHF0U7uH2huxE/quXrdYxcfusahH6z/kFfcV
0anBWd2FyclhfGogrG8jPyg6XiHpVqM273lkL7F9Il5NPqb5Nr70jDb3zRNYmIoN
krQ0QUSTwrcU+RFUqrr+vIsjCtbHOS/FCqzon5Do1YMFQvaDiYa2KBqxmIv/w5rF
wz1CBDzdIXagheacUQqzP7IkkPFVs1ZV+o7opveHtGzmFW8HZVDkpg1upcUWZN7A
UXiIY1nYL4mNtTYund5WYTatB+1PrLlu5muFp++awRgInDEr/RDt+ZA9VKwER9fi
HFZoZImopxLp5ZWxNRpQH2SxRBhEc+PVIgV0M0Tt64k53QAQkWjOvgg3vlP1gdOT
ehNAxNbBzl1IpFzU89N5XEM4YO285oIIBpu1QGheNmwrVoRC5uiGTzkhgKVLbpii
Ue6+6yJtMzouLxIisGQbZNem8uf1YbVApxyYEuKnEogExaB/YDwXqDvClvqy/RZo
wISo7FJo8Vj3omly+W5MsorTT2FXYVO2Ziupe9EPguIf/YKiTTAHmWJjbMTw1Gy6
Q1yuph43PJYzKBZQd3OsB62EEkjVn4A4LBW1CXLmlCVtg7WjeAv4AAeKFjzFtuiG
ycWuUN29Wu4f3/ZMZpo4BKNVcgsiOi3xrbEW/fc614cdVIig6GV73Ugy/qYgru/a
atd33eAHC7YaAd+khZq2mLc31gUsoLpbFlHQtKlVxWVRQv2XcThMsdZklj8caEr/
yG4/LJADqdDnFoH7zEpDbLMNvwZfsZv6IFDtlnYCAqscdpB4p7bIcj4AFbf1XDO6
BJy+ermxzj3iyr37x2bJ1KJln8MSm7hOr2yWFJNOKYeMUyHwp90OJkL69vOtMRCQ
dMv3iEuPTkYJzkRv8gR9kxUboHZ3rCXdCP7p5UCg/P4V8Er+BUpkbBSpRYPifUSX
uNSIkfH6EgWJuDkYT2WHkR/shQpw9GGGx6rwjpnrpzQWnkkP+s2a8TTZakJnReyk
cBu1c7aGy+FhMq1w+XqaZ01R+PWsgnNPciN5Bg/sNn73Yv08uCXvT9DnT/p6dLud
HjbXT3q9kPWJmomF5t7rSCS4tYsR8EeuJuP5TRytA+RtKeDifGtNgliE3WK61ToE
+3vjcu5YgKgtNRES8MPlSVEOOFRwz/KXwFMe6j0+l63rneYMDQ5Yf2Cuo70oHN4v
3P0hHnQy5V3ZWB4G2QjeNkki9VZ0jLIWF6Vtc4FB9bvDhSCIx6trKj7ieA25hj3R
Ryywt2/d5CWMa0QDWmESTEpRyuQx7Cb+GaJXwi2bbTgTmPW+ZiOcVwtOpzI6z5Wg
6cjTAMWUmop3KpIyllAyfIryhkj+6oA/DCTUeh3lab/tThV+59/UF4kqLgsSjvg4
Of/h3DX3K/oGZVIfvkSjUTb3vwIM9RrkASOx8Ephc64BbHQ5lYGZj09VqgWDZmp8
EcdHE1ZuG10hPOfgGpql1GPuluUIKrDL5bNwwiP2o9X49QEYGM2LAg2P7KV6TW5C
lg7DOdsrt4jmaVjGPkm15hPZmYqnOHESLwxZQl+ejNI/gWzOsqCR4TPEYtRXLu+b
uMUWd0/eRwOBk2Yv/0jePprdwJNaDSjCg7OCCPiPkatGFEvDWlSWjyxeVDSqkcEB
YIi7nbg4bARFVShkIElVYnXwQtPUZFUueNCbZMs4dgR4EvjvgqCfEkFJZTaDMxoT
jDSPd052XUdCpZfO8pifQCbngLDJKdvjPRORJR+AiY/rWUCT1g2ZQBWdTcMAY9Dn
g+2RPI/SLY8BvTRPIu5s8yUZ2Uj9YNIKGRVw4lajvNp6QDYIKZ12hWVRfom5PmMo
yRi3CcPHue451akLsV0/o89uW0CzyI7hlpSdro1YGDXK3arffHyKRkvIuXLXLsX2
jaLZGCFJrRQOvhZhKgmsPrWM0oDtg/33e7lQDnUO6urUM24BGJgXCySYNZbIy9NZ
nhQLpQU/k+fVY8ieZjCVYDcjp0rbsyMZUHijanAPSRfp7buRtO56msgTd31Xz8fo
Lpv4h+UeePRJBhn//SvE7Av+MRHGjR23qlEO5YW386RjkgeJonXceD3/kLThoRgz
4RDlnMg45//BIenQhdjk22L07KhoKydc4Dc7BBNRNWShV3k7dc3FPYkvujgOzjmr
xqlPoLPfJq8/NcTpLvzXdfQ+8hOmqhyON8Vy6B3xniKviO0bG6ctiRQJvCv5m10Q
Uka+ETsIAqXMCTnX3nJw4IYKmSLz0tqUzxF2G3TUh68blalgNmL8bONgR1imOxmT
V2QRnUneLOx+/Q8SREMo6vtrY8I4Vz1hK/2T36y0390dyTAiDGtGcQnYETsph4pp
GC8aGZFbneX2QCcZsSRNsNr9OCpk/5IjyVzMQWzgH8LPbn4Q2ZOHXvn8iyfcqQOd
Tqc9JiEStm13ENzrNgkambDNhDTuo2gt8ToBco6zvQSsl66ALWngIVnFZHmIjPUi
ipwTt3gsb6ZobfbZe0PezVELghVmIy+NStW03wrx4qPHYiqItDi9/GIQX2dVO6FB
NDw1V3UPZoErwsfapdvefk7ph/Cfz2EtoJqLDqcTru6qXUxZ9RgEI/zfVxzv80ux
4GAPO3CcERGaYGs6CfEFAzrgpQem91AeNA/hDeaVTcgjjBoPITel5GBWxi8Xv3Q+
g0OJrdyLDFYC9S7FNRqNB5fY/deNmytYjuOeM85KH+ZIDbeYyzjEnzFA84Mk0q8p
ahAaFlcszRXALkzGTl3BtCwF4CxQgNqPazJvNQ3nz2ImOxTQ4JDIrfLejP8HHTdq
WHU2w0U1OuSG/mTb9hTFvHhurNQMYXjKn11pi0RyFkl1Pt1SJvERYs9Zgdd17mM9
uB2W3jkHsZ6bcjaJLsCMl0aRCRNEO7Iqi/4LJMCYAUXuFtE+cuzx8iTtD8OX8azD
RhK4TajI7Uz/6OfYNQoRDCSKA2K4vgAuflovs5iQQi7GGP6/ljVpItvLoXCUZTPZ
UedW/M4UVL4CSIDTRIkDiuIAPGcRLzYrFyCT0H0BlKhDiYqOByIP8WehbrAg93cP
DjFKB8UpV6BcjJiLegfG69RKVawUXPMhqgNwi08RcjSG85+AXbNXJ5tfj9ekS5rX
ai4KSevXKE7Qeb+cEoDTbubPmjFuMgliqpidrVyvTFv2szALv5nFClnaU9YFIOOq
B+IuFSYTG4RXg5p+fi/PGuKGQE+phAi8lcybxUJhwU4fW1FV1WqyxrNZrLiR1XTw
ixaI4+6iiGFWy2u5oJj/1BYTrg3Bh21rHsisuFTv3XjAOyt29fJkhBKgcuMUS4oK
F0nhr3QiImRJVUHS8BhtX9R+v20kSksFOH4Yp6KaUk6eHHNaevb9lvIkcZACt3n/
BbJvSxgKSBGARsMKYc19BfwO8pZEvU8esGCqUI8iunH4wcBRmv95aYbv94RARZkZ
viMAiP8S4Wzjr42oykVBUuaLsg0aLQB/0sCb60w5HgT6/hf9nn560l228t7XKRQQ
pxoA9o2CQh4RbRusjxbwTfGUxRmI9yFYdUGlDBNyEBKzsRvNTPv5Ly/tYmA3J2H2
4jHVmvo0joljR0VrPmTIj5YaJJnPFG9N7iC2R3XszXjKshzV3cCirEXsVGHIbgxN
Ov3N/0GeOK95EJDl9XDrQRgHmlN3z6ZShRXgdP9uhDqKwYm7i+BJAgZSqKgddaCw
faIGFJsIdwPFUWfI/UoXQrRZWMc1APmx0tCNvfTTtsmU+srAHmxUTXmDEz2yh7RY
CBXY+Ncze7586WkTL6ciLc27ZwSjNzOPmhGfVCq0XIQhYYnUWC+ATcykrqINZhR+
0a49zMc5j0hxfbsQK8Mq5pcuf7sigdKsUOmneghU/LvAUFp5PfVEWXhRsAM3eX0o
8rcVCBuB93aS8YKG9/5027x3oD1e26IHU8HLJ6zHTcW/0fLCEkYeDJzpOPya8kpX
idbgnEAuUP4riLtwPftl73zRwD3eE/3GfVxhOfjkF4TnrtG8ZJSSPgau04ngx6hX
WVkDV6L4ZyBmOIX+mL2D3kf131PZLT6sqErNgOMXoXSHLnrhcBkdqz+jmw7pMYVA
RzxKCWAV9oiG9y7Ss5p4KSQD9Kf4I37aAJ5vNIyVT1Ym81r1D4+66NtxT5GFnYwa
nFiXewuIhAnszt5ijkb08nNFYumv+avri0YhyeL7B5yB1OGUOVzVvG10+GsFWBpM
iBmMekOmj591eZUorRU4+HVPijol4OfEjGZbocry6mVgogQ8JIMKVQ5xZAx5qEo4
G+YD4f5bc4pSkufk9ILhlu3hwiO7FI6qbqdRJq6QDCubGVJbD9e6AsbfNgXN77tk
1C509meumgjy8LEtDYqmk7zNiZ/zylO0YYsI7x/n6eM1AiSCWe73o4Sf69/NCZ8f
ZQ6DGo8+c3NMRzR1Tfl7+JEimNG8pA4i2MaIOnt5bHwOqqCb3/QqbZav5WoxU9zb
ko5fBN24rns+SrZdw/uxJvzwZrnDqaTe/zj/9rhfzmsidy72zGZX2pxJLIlGMq6Z
IwrO3SqXXa+bqhBuAZv2AU9Jw3hfE8xfAHOauxgUPam5cBxJNzL5DI1IEpzptpSz
1RU+8GvQQE3tEULjKAI+TNTtpmnE8KEScR01HiSVfUV1FMNJoLOYWnve/xreZ1af
Dt0N2NenZiUwlvocFzU/dtvjlO9b63GDT96TGQGzoYhC7gt+PnhjEIH+8HmVHHsp
1uepsxwUh4fFxJConVF990CMOt52qkMeGSoZ8tnSD9uP93E//O5yc2lXr781Emy0
uInOZJcx6rvw7uT6INoJmfui2IgrzVyKrNrZFu+R+yAV0ve+mosorl57kLSdKino
KUnONrO5+M9P2RzDm5f+olSWiI1TIfBjX/RLPWuu3dNkxRdW2CRncSmZ8UVzsdXM
UNcpHOJvg8q38C/X7WHjuf/Q3rVW65JVjO3fTKEIKy+kifHuuqO6zkKQo0roseNW
RhxTcl+iKVGwAvlcbdzBmj03yT0wBSCW0h8+5PSkHV3foa3NsJFpAsDpyIDUSoqk
nJlvQ8/cOFcTwCRXYtH2oJEyVUOOF+PNzP7JGJdTHrxvVgjRkqYUf6bBJKygxlfy
Os7TB+iJuGLNUREIi5l3c+WjWKV8MyUlRCNpeEHkRyik1i9QZII1PYs6UeUICNUt
O+nkZZBg4qUIbrR3aD8fnzrmstdYsXiKi4BsoUOAnBBfuQYwtE42GGK9tryxvUc9
YCP6766PHQLAjJuhvIASp8/hkohXI71uhKDAMy0PoGugonosyjRUm+Dwt7RvxtbA
ATomt7RDutqzSNIhQvCOnwWg1DWH0lEHZE+tNFEzCYwTf0jke7utDIdLJesjlxOh
e/OQ+/0cLB4FmzV+I8NqilgJivmB3wrOZsYrucEXVDWY8YjTbifnTgOUGW3Bun3v
BsjCgWX0ED7CQP/9INutLjxegHlG4xet3b7s0RjaqZ7Bzn/h3fAoRYna/cMf1KMI
WX2xxFbz34E/IyfnX84Zry7HGJ8WQGHRHlWxK8HOgN8vI3TXwXb8e7KO91Inw6Fi
MP7mbXGfyML/V1BiiZSn29Jb0G2K1uWEoq+1MHXefgt5lcnRx1AmBM9mNR7pAh7b
CZxUdx9nMLeiBft6A5YjCctN65q+n6y4ihDJ3nKNa8SfahhIcSjdl2odgmcEKuOz
mnwIlMiE7WX59wBHxucYDhMpYC2UXqUCbQur+ck7rOZuC89hED161ADpcG+oPT1I
zHa63Jc/kIClPeo3GnA6gca3f9tAXmm6I9dHS9ts9fq56sVvlnm8rImPe7OEuT1V
jUdYR0gN1pYhDKd6FxzWLUauM55o15E8K78JMQPbZVuMBatM/DDOVKfiJuc7DEi8
smHjZlRsRwHjkIEngV1vTaxTRWOTSAniVNaz/fRohRgdHissePRCLi+uoaI1cpMS
5Q1cprhNKOJaPpLIKh7mS189bpEDiUsqlauER5x0bYx7Y8Y2Bd/JuqCsk4p/6L1k
Dt2BHMt4UPk9LgnzO3/rhFA1o2iDc8a6puo5X8C4TKV4IELCxf/uzz1ysHUSQn/G
wX+Gh50rJIG+0zxIyfyRFNRoDJRTG4HTaSIbIEYdVgKG20zxTXIQf0/vUdgpqbjd
jt73jH4QdYkkzBjyaT8KNpNbQcjM7P2ZuvycsiDhRq/LQ/oq/D1bwgru0DvJpPl7
ITm7/65K83sOCPygqMLp16bgPhCZSrdF14hlfmM6qa7ShOebUQWhy2Sg8UPySyFC
lwUiIe0qhre5GSsdNUhxbWwb9FFPDpd3yvcGj7pEZCpu3bs2nNSjzlUEnQbNpKYE
gjLSSzYDbesICwFDLPMXyO73s1WKlZkIuWEZnXcmQ2Sb71PvP9TWW7nWwQoFWoTG
oFfNNn08QGnOOXsDgBRkSZl52sEZmJ9SkQp78Pz9bQ+5X98Q963Hu4ktIc1jTQ+l
t8PdihLT4B4884QI5zCUKY79UdETdhsab/gpvyWEW/4UKr61GrsTbLUCO6QgHD4W
z5XbZYFakPyVF4kym8593RAumK31u2UiQWD+YKgwVS4/VDe5GiOy/X+0gM1v+rEY
4QzMEUlQUH1EYFiimyGr7JJ4bFopz/YZ2uM9XOyE7Nkp3H/Nx5GP5vBZKT9DinMq
1eHej5xcbMzIHWrEIxcIJfk3f7nOZMgko7ltYMKzvel/JLFmhj6J+JRYsTZATDcq
GtBRBn4uwXw9FHuFUWU3rw1pYip19pqRqRGCtdeMB8QAudWWoIrv6M7kIJnwaI6n
UrAUjqwOt08/VzhSXWMWwIP9khA36hP1YEdsT71z0XGsb+GwpMnuWSI3NFHRy43g
Z9yaIlUUE/eDIJE4UfZJiRY3FPDsLHChJ/6vZ6lI3nNM7nARN2NirDbgqjw2Ry/q
+qnKRxtkj5A6+Gt9ECpxyf0qoA3yEs55pTqoWH5n/pMXbFESiHndcDNiUJHgXze+
Zea1Gd1kXCIVsXFoejfgzOTSdT9AihntGVma0RN5EvGRLFmxVTVP5lXGhCDSt2XO
PEYqPUFdfs5WMeL96ydzcN5ZTt8Ll5KP4mT2PObcuiLYn1eTuL9/rYgv6fOq9GgB
OV9qEGdga4NoDzVF8MnQ0PnLEPCoCm4RvzaQjzNLC6EpByaGH9QTTLiPUGpztQmF
agmBtM+p5Zw7G6LxIkR+bQ8oA8MvRT6F/SBXXmKDRevkWWFlUt4BJtWmAOJAVQpe
9ics90v5Wk7B+f0wj8Pmm5JGJbXBkrKFnVZeLIhU0AuRv3CK6+HKngObf7C+MPh6
CR9OKQ6TDc706CG66u27sr3tyniOZCntiKCT+XJUzfYXD3s0mTPOcxqjTHKdqj/1
FrgV9md7qJUppX/QQaVZr+cCWG2T4ppnCCNWMwcipHHqDUt6akQLxkAtT5GTXqNu
FGpNZffPJfCIIWUJl0nezahMimcggE/ALQfUCvegs4JS5EjX3KmsvcjD4udfnmIm
VVQ8awyyRQ+6TJGBECJ9fOLOC0lFchbxHh9hzA/omKYasduH/2+Z59xEt/9dMAmu
7IYpJhCA+XXvogAfy8IqlXO53N3wswfGpm0M2ZQ6ClZ3p8Ur1bmR0g2wm/GunsBL
wC64ZVtvRio88AQlza3m+FRiTQkMETbtduGwah5+qA+ukKr8rp76ftO/8KFyCJVd
yNYcgw+uErGOnl0wkD+y0Q++k3Vpd4jbawemHIVfsP4gCozDfKiaPJjCoGDrovjK
vFmbZWeiALIkMLKE7pFu+7N98dPQLD6ANHxgX1ZjhejaeRYTlGX+OjaPpOvl1ZNu
C2gF20ge0EBhcmih5jbLxbJJtGFM5PJt0igYf1ZIG8XXsZSdDkSYC7nNW2Tqu+Uo
1Q5vNlTKO9h8/l1jRepQBYlTTOQA8EGzicD8+NY2w7rjuD0/d0S82k/l4s2vx+kv
KImXwwzP1WP9NySoTIRIIxJjYPoIRQtViXLLFSxYUDa4eOQbd+ZYRsTSTtAlLcVE
mbyD3RdJ+4UqSetB3GsJBzbSTik4t6HJAqm6frhYCYj9iWSbwqt7B+Sk0C7aE5vc
Ac8H2dS/m/lfQyR6koIeW9NmiGSYWnVe5jBlcQvCHJxO/DZk0QHMjBIl6gnrzsSU
iDD/ItoqLY7XTbJRvNJ62rpxiYtnRatmMPyrGC30riqvl/IroZFnLUFfRlElvdWd
Eaj8wVLNis+5C/i2nQhg3PfYF289GMZ27GVmsLC6ura8XLLe6SjAaTuyAOJAovEJ
eybK5vKAlWORBQA034W+paei4aO2XhIKmm6N9l6H5cNVsDXoW69PfJBeoRXdNZAr
3XeJsBdHecLh3Lr07Lfhs/UX5AOmdeTRTbUvtJSLOrg6Lxw5b3pXoOgAPjCcmrRs
7CvIgAtY5w9I2kErzqszH9lgL+UDmirHgyJliiALssWdWvRLQ2XC6aqTdW8wI/vJ
k4zgUn8oHVF8DhISR+bhCd/+tZISeop/xNYMGWdzRMWMf5q2Mvabq5pZeCZtf15l
mTr0VCGXahBRgrspS8wuZFA6UQCuJxefvnbZqFxk3Nw+qszJ82pMuZlpp9wlWtN8
H3hJTVJYk6GfSDN7LLGF3kmXRnoMR85o/lAlBby2w0Rym134WLz/s5oKZ93Xfkb/
rTYNuRLzRE2n9zGu2XqK1KHAfLLNSNTGw+Xdgkx0QgJEwxGS3LA3CfyVgpl518iW
uR3U8ZbbhOutOxwBA2Gl6FY06r5Mt13QPd7MN5gBob0vbHVNgUZfj+qqKvrGu8Lu
Le66AxDObyE5S1rKfvuDB7W4FlY41f7gGxrunqyEWrTbsd1MAdD/qEEm0Ax0V71/
T4aZks79BG2aBQQ9VkBbEC4WVoh0+n9c0l4PacEQruXAuajowq1ZWian0RnFkljg
LSm4/WPpifveM7FS0uFTyrdm8KTB35Fvw3zkAyzvZ613UHPCK6ZIf8jIyeJjdWRU
Hdxi/3Rk76zqjwtH5fpzVdehmdUt9cxo7kzTvye3R3D5BljFoxE5Df1VCDEDboBg
fuQk57ro6G/RuMZ6zR6vfJc/uXPzaCAA6XZYVEsAhdBD2mTjYKAJLP8zVUq3ScfB
1An3y18JfEQHUWWNXOmnCWfNOGtz924unYuz6ebwLjU6PHbzBEdhv2BR7WIHQ2N9
1pzRtiyuZYvlKNqVvzcwqA4Dq5n/bjZP2LOqJnNSpeY4ahYBD1cwH7rta9JXSjGw
m6m2Y3rqKCvpLEGfR1Se7U7vgi7qlTtlswzw3jdEsM5ughjRdrCnxT0iVIQ/r6ng
atlaHjvRqJITC2vItH8otJJW+gXlwKMmR6zEoo99QHSew47ydWngupLgdeyAYUgl
h+t9h2dR32ioraSwMa32GZuhksmYfBneapfRyqMVT9uizBDvi+NAPuD2pnyKX34+
WAta5DT2VsSDRtzsW3/3A+y8HBKUWhc3aZ5e7KSlWz0ciI84Yt+jjUry71N9agF2
hCiiQ632XieGCEx8IWw7+Cmbf/08JRQsPMFO42aVqR+WDdWO+8Txl0RywFNLyXIT
HBBQ8F2fphclfr2PfYWBsiNSNcw0um4sKt3ToOyCdQd9oVM5IS0SLxkDQUMh/3gC
HhOLSDTI+6eTxHWd8sgE/8F7ub828vWA30Cz22le+vAXp702pQoRrmlnPRiqJBrS
+rGfi0K4MnU3B4aDZig38edNQlXOokh2otElIes6ex50H1YgKg64xsVyiAYRBWSE
81ya/sUQERouEfSRwjEin+wH0LgZ6vs1wbvzeA1Z23/1+3PdPF6xNeBELgwgN3Ut
6EsrTxq1cKyx7+okbCfsn5h7S6LYbHiurL7Drim+JeI=
`protect END_PROTECTED
