`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1aJV+o5EkDm8Zrc0haE3ZMA39hBDGen09+WNU+vmQmiDTs/hR1Qgn5hsG4lVcq5h
kTMRr4eplQfr4xe5DpZ7Fv8XVfx02G3FPkjzSDpcIHLLs2WIz/LH31GvPaCnVzen
mrkFkC5UCqOC4/KLDYqyt94BLNqBh0CwaYW2bGcK+Vcnk6BSA0eFfq+rYvd1iT0n
r8C4KigYHkI3sQLK5whiEdyUHQTum6G8us7I/qIWDKzKAjiwQVI92J2sqwFcZlfL
w/amjof5ucu8DX6gTmZbIHSZ0lEM5FKEybcoVsOWR3SNT1Mnx1zoSLOpmuAsXaJQ
pDrnUANt6Nwqf53OQ1SQEEOBcQTRsON2QOk7Dzn0fZmb1pZe8XgqWNYxHYSYN9wH
17RRwIFVc5X1FOM2Qbp1UuBpNHEU/0QhY/zaAws6jxyQwTE90K6RAYNOaMCaZq/X
Mby79318XtP4U+YuL+9MLp9Z9/HkmdzKKRs+RP0ussmWxk7u59Dm+4rBAZmId/VT
XDDJ21NrDlOBx3Wh1HYo9Dz4CYwBWp+QiYCb2cmMCDIWylHhfmTYzitSM5IVGeZN
vaf/uY60Uesp8dwMtmf/GcvuqJHpFbQU6KC1WsJpabUyOUovaXrTd6rGCLUyuvbT
V333z5nTtzjik8q/ukBxAG0IidCzbF5zoUNe4kOpduHMai4mSEJVitQ8ZKQB5fZs
HRF3qPxYHHbZPjBR9Yb04JnUekeCOwVm1WL89D3w29snas13Xyou9hTLUPZfQ/jB
Z8ExZiZPbuf4bWZOP+iF+g/AAOTf+FhUPnn59s8psAsgSor0Fx2mwRQVbk/+QybT
PRgKnOGBFcwqBWhx/M6PAfKZcyBApjr/M8TuMdl3+XBJrnxheCzngGDVTVlTQ+KF
+xyj3UPdzPZ2KiOtz1FNBFSMuOBurDJzaLm8tSAF19liHfKOCbiDVIlAlRUjd7oX
Io2nPo315i/+42jCwqLknM4kuQpScfczwtwAI+smSMm04b/bvNsKQb96dPYrqLz1
ZffDGvJRTioS2gvzq5Mp0mrFM3Z+oGESDdIGYfd+FHdpZ/vTShU6qVsc0p/ME7k2
MKHpXdtiRJag8/aWYHFQH+E6C9vZxOKNabPbV1G/m+Say4909Uz72qW10laVEoB/
z3Rr83aNOuzNrjY++EKuvvCZOKhJo41hGorblep3L/v8WJwbnUD7AI2JVv9MiQYL
D3O1OrXlWk2mwJipZp6Mo+d54wH/J88I2qHWd21OgXRaB8cvXyHVrh9R73VNDZfg
QbgM381SbBVHvMtJ5mvrZ6g9PPnTRKuxkQEzpxRNFcR/SiKYeALSEPPyfKv7M+8+
+FBG+3zyDuENOwnGJDXtbqlVcsJ6/rDRGe+InNJnEJPOZKFohM7hPcp5YfGsj8gC
Kk3EgNau7k1owPLUyTBMLJu1NIdqCxMKAF/6rTLWNoxqVzx0m0kV2jByfnI1Jd2l
KC+TyxG3USpO0BoJHp4hPyORJVsVZdrnzdHrmjf5d1tHLNntbeG0KEIB55MK8uDs
0fUAAhgMSZumXJi3LL5r3PRbUmdTBeKHa1NBQMtauybT5bcJHE4hHCoZ+g7lrXQS
5xb60xC+zKi0l93YFQAjrvshAiMTkkyBmuPt7AFnET+sTTsAVPDzEBV/7HJV77lT
D+zBsnJVDFI/pp52fTMSjgdPVFqPcAnPod/nu7iPhP/MzhvzjZoVenfnoDA8CI2z
FUm0yVCCnZhUJXeMCxepjSIVP9oirsPyr2GOrK2hvS4dMOt30tJ+NtmYvCV1VM6S
Ra1d+lQk3IdhKRMRDPgVoYJyfZO4mTRwYu9M89SeNEhm7pfitaZxPeg1+guCejm4
hYoMu9q4NrL9Kr28aF0RTBLxJf+IGpv2IqEZ7A7Y+HGDdVRctDR7cRvacPwfbgYQ
eCLS1wI0Xrlxiw+ip7LLNN/aIJ5QNXLgKSgHAypi/6ZZSj3OWtZUH4PZKwMdJycr
q+mNwgvU/nQn4er7eFMu+CjDaxDqH/EFymulE17ASb/panstvce9hfKpk9vXMhYI
poHnSY11wkNrr8OegBgdOIAb9oKvvqXCNubJyWIrUMs2ZiAETuIYKRMrTfJaBqnF
drBumwqDz9ZGJlxofUiDtICZMt5ykDzX3JqWT+M+Aql3MtJCdIbmVKIMpfvPcpIm
d9UccL8YVjJue5K3lRrpKG6iQJZSNgeCPj0YHX9NyNHsfQzm9ReXNIwLvc9Bd+NZ
3VMHyvJ150oPFIotBgSv3U5MR9pdxCUSk0mbVlZpXvrBjXSQrTRvsPE8U4/Z5uEh
7WwAl75yb/8kO6q8ETOj4PuOl590v+JkXjcvL9Gz3+9Tv1oct8rc/8b9ECGnzqzk
zePG611YjoHw9kO+Vm/qbLitzuwGmwlw4nV1/1sanrZu2mp4FzAo+EVreYvYH9hV
KiPGl4RUwGk3OPSt/8w+YbLKIknICLvjL/cJ5ppn2athJVCUZiNPQcBJMsdcVtT4
M63EKNu1lnNqDtlBeA/r/a0yBWqwbFit+VvJA92EgiEVYF+KtvCaIfnxeRy5Qcb4
xtJDPfOVY6o6l2kWYq/v+qA4RpCTbJLdAUSmCccF5t4cyw+5V7q1js1sDwA9hYBV
o7mqBFiU5aoaw5IyGViN1k/DE8AidmXTbMN8knUP+Q9g+WJJTW0xEKXrjrhuHO7z
4Vqqhmrdb1ySQRfnFWCVMjJpihWWRBBFmnYE9O/ibUKUH8Qdzdt4dn+EqMLIy1/i
y8GqW56/v+OMpR0Rg1nSwOY2zuXSXsUYRwnYXoiUTqd8nCewAo/Suclsc658aRYX
bMDvuBJZ9ZTiCxdjrTGZNoU1k04/uSqhy6ba6GSVCQ144IbinvIJe5vYPW7dtHTZ
RiHrr4j50AdmOx9Xk5qZ/5t3yoL5ZcBzt/MOovqjqpovN9+YM1M4TAKQGjZyNFdb
ChPFAnqodLlCTrYd1dxNEhbmifh66MBJcN4DlLrIm32yfEoLkGOxk8tJyMt15r+3
6WUtJT73Igdtc/CL/xCo7XBP42G7NLZu1iYpJZqhqoA9PH1PCkNysQLbDsKLxR4k
Yzi0pM71z8R260rBlFSRPdStXJCNfUcpYzwP8sRrCxn6pYyN8oplXrK1ZPU9pUPh
RPnh53gr2tb2RHCs2FpQo4qNG9cUtwLetGjWkR7rVdkO1TsnePcZ6rWk9WvYhwd6
is3E6cMOabxKFXmLjKW29+i9/rwl8+f7z8ABJd42ynNG/AihgQfMvn+wTPnUT25J
KvbMvwGSJ5EOhdfuahlBijoifnzydQBUog+rAChfcQ2f9g1TzMzlDKerSgGTLIme
c903+RcLGZXVmyIiRQ60d+YuPoxklMBiUdWj7oz7QQE6YWX92aGXFUbgzQcZwLsA
FwoOtQu+TnU4iHd6IgAyOG4wz1A6WvDJeE8Zi9CNJAGxWdjLvu4rnpmS9q7416N9
YWddC6pG3SysaL80/mAJf6cdUWilTwPlydmBA9K18keeWO2GiONwUnwCpKfMij9c
KfLR9vVBMt89xtWb7AHfVaarTKFILbviJgyzVgzbtcSXTV0Ga8U6aPz2z09xKj9+
NS/1WyaoFJ6SP6KZd8CmvzcRY5PXbNGDD68Wll4UBAmV5z6Bwi3arpCTIYBEdbtF
0i/4VBNjrHQEnRCieFM4A64lGIY+k0BJMNRSUwsBW9sz/i3TuuxZCVAgq+qapXsG
xFaOALmOzfhOXlDd04o7i8Vs3AF1c2k3I/FnD2r+nPX767UFrk9bwcZVSTqFngpE
XDeuJHDdnCOvhLUeSLmzzLdKqFZPszBdAK3W53Sgek652F4N8Ig40aue1zOjbyXW
i69c0W3bJjHSDaTa7qD1at56rZUmAbcBLOSO9G37L2RC44/LKnUC8Cy3WtX9PZoa
qbb8FjyvUnJdRiBcqfPFRJECZ05dDHbHpht2lVG8wXDT9ftlFURONYj+ZOzQnpTT
CBynnh99CTiOlWLPrD2+mMyhAeljAzebW8QAIkGDX+nxjv4pqSqvxZlekyzUAX4Z
ylQ43RjA1zzANp0GLV/nXSGZdp2wDjbEztly6OZCO48zK+Kn4T7JNaEFIoxtu+L8
GeDVGx++N63W3MYCvJLWrAYgGhWLKwt7aj0Ir4yYpd0gsKeJQAPkYXnVc+AvUuen
uUIBKJQ8zxTqILDsjtaenlzrAI5+xgsertRXp0JUMRitYXvXMouESI98iHXwcLvp
EWwJ9U1ysT4Yaqjo0VcHnEC/N2YRZdW2GW3qHE1RpSW9IG5fwqhKweUKEJbXxazD
1njiNWOmt3beck+cYu0g0VKfSqwKTfng52u9KLGWHYazizjd21hIoUWGXXq9F0OX
dlBFyAx72HjZLHw52WPZoDENwUn1Q1hReZtZ/QOPwJgj4iXB5/+6k4VNZ5cMHiiI
GV1nntW2vMv4fFA/+1l1iaR5hJeKnRJE6bS6kqGQxUKs8bp3221CnGWB9B+URnO4
E0fbV6YIlC5qxlpgbJcbHElH024xob1aGDLZhOCwOzedgyO9peQmsntBz4U+4xB8
T7NMoNvW3FPo0LPZBxo3eVzM1VUWUwvoIKWv5LPiZZo2LLyaSKZHpRpWNjtnGcCv
MkA4XsVBhDQxTaoJr0fqgJAAfsGyazBrEjMox0NCDr7GGI17UTrEx4oBQieQZy94
ZgI43E2T1wrZ8KIu6ZLTSbmtkJ7B2JipSLUxPVK1WXXPhdz6eTJmCIz+mrD3BHHd
VKorSQsDMRdwFGm5yUDENEnwNVSV+7JvAv1iOxriMw36IljPUI0+FB0gjKMeY3il
LBxo//+r8Dqy2Qr8EKUiSD34FGpK/JIQ+GzRpFMPHZzib7JBh9Ph46GUEA+0ofaW
NIEK6xGidd+03nzyHPNhR6aMYiOHqABZGqWrX5iBDvd/zAsB/ckHI16C9+VfC/1D
cItQHpyZ6hl7JH5rtBqIAgZ89S6V8kFiMCcRBWiAAEpljtPmUBsdAE7QPcyqcSeY
QSz515cJaGC4Q+MLfBVDlG5g4iyCE5d871W7CafdDn30gU5kMmjGzmNPi0fSRpfs
6Jd1pAQ5JAU2nxC7yuGgJXKytrK6MF44IZFnwZ/xTkA3jnPP9VRi384VgwksY8dh
fcGFnXRyoxN4MZC75lypvyDPBJGHcyRnDuD25YGvipcNSZDxyJ+zl5Nlop9Wt3hu
NrhPQXj7FPaf7IRPDJRFhvK0mOTClQv4wbjOho6BTQVQXQT0RXS5LKvCaAaiscFd
gq6hZgQeAbtBGL163S1xCI3hPKAxi2yKPH4znTi4+/6jk9wFHnAL0PuxB7yS3Tyg
VTC7njN8YNSgS3vfXPMI1aNNMGVbWcIxq0cVapf84VztEq7cRv3D7oAk4sglXTs0
bVZ4kjSbfCPRA3uJbKq3E0NLoDE79+AfKphOl/vCTNnCH3FOgg0CHI21NqafrQJB
9ETHIuvlmWkpPhN7PNz1xXaHNslByqeK+wS7E2+f1YTt2PKzDFhmb8WQy3KZLj3i
cDOG7WZvAEgBtq8viWvCkue7hqXS7UxPWYM3AQyDy94ZORgYBmic7polAnnUkZY3
GBXKvIz17XZuPbN2zdmJB1w6E8ym9AOFmxFh7KymamjnGdA9nt1Kc1aqMuzmHGer
BJilkFBDCkDMirsZe+m6emvKd0MfdeQPqUZAQ4LgeyRc9G4CaEtJyCKv8LmobDhs
`protect END_PROTECTED
