`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6b4eLmv5BXYGmi4f6TJDKte55OCPuctOSI4Wuoc5+pmCSAfNZi33Y+hmMGpkMU+
MOS6OgNbkFMDDy6qK37akKtF/TgIvYzNhEMw0My21C52wJoD3waazQ4LOdmBcDap
F+LlUkzIQEtF5PIk1gXQTXIuy7s6Bs87pJqm0G3WZ2Rh9c/hgkRo/zKl3cWhg9gm
yosAHcfkNCNEeyb8ba/MdHM/ZOP4llBOTGK1/Nzw+vWsqsGjZ1MM49YHt2q7QR3L
YNVqaO++OM0SVuGXo/jlhybSQqxXq4CRT7U3o9YzImea6L5T9NX0vXONAB4qeroB
PKRkkzCUphb5CNgwqg3eir+QUUleWwic6TDu4H5T7DQtI2Mw7lMlXCBH2RZTEODs
Hz7SdwBKgs1WB50D3rpmkB9Cg1+wQ3M//DKVDVofQQ1tLaGBSWFqk93vOOV7KAC+
CR1rlI2+cFZMP+ij15gXHLCFSD9p7HCqPRxBrNL24WaEkeo0yFVe5yWv1b12fWFW
zqtVTx7nAUAeJh4+0RVxV7r2Y4ejF21/bucknI8GK+pxl+e6EYRII4z1+KU5i2Rh
TdWNsrVeu6dQ/4hkEfFeantOtHHi9WDWyLArZmrAnIHY8i6Qdn1mkNP73h7UAN9F
cvH4i5Kj9XLLZoynKFU0cGaDHH4nT1UYADMl5epAxdL+TVFE4MFH9A+mINmFH+9v
MXnNRIPhJQW3BKCzW1S2y3f4sM/1uHW+EhUhX3KDx8e6tmDbza2DYpU+RuM3UoYz
VA23/T7KQRZXZPdJzHuQcAibii8k/MRsCru4b0Iq2FYBLaABo8XrpVIJX6BYw5Ag
q3JfJ3AvObi0S2ad+UswbtZWy0zFKoqy4+MxHgJB8Sfk7cfKI41Vk9ZEPUP3Hlgp
BU1wJFzuEWlOv5ZPZbXK3dNyjxQdRkCw4uee8rqEIEFYXjBBzS3cE1Iub/b2rXeV
Jajjy3XOBGmTm8SQsZ+drxH/i8DrNBFPBcZjMbodXG9DshSFZbJGUfj6FcbZ0gkj
yuiQr+sebCTOqNV8j0/Mu0e1fvIRYQpyH7ZtdqXt2DrEn60sQvDTvG4YcwnZXBtD
TXYZuT82ufJfxWvvVZYSO9dlpik+yKG+hMGA2fphI1ETIKN4RYHSNNfOXHcPWXK+
gVZuMHd2TaWCXSRumk6M5RyK1saYuKPFgHwRIJ92PstkgEagOqJIoAQphSSHbSd+
t3lvF09+M0XW8zzOmkYmx3LdtMPipnBqvr9IDVY0WBKFYI346fx0wzvUWnptIkXS
/R0oJsRBLASgukg87S41b1dQd3SyhtwUj/7U+t5Go/m2cdyvGQTs3yj49AN+IJKQ
DconpcB0rUnmOB759ZNHjpamC7wp6p6lhil8QstjQAUtRto0Ao76eeYE97yyhFr8
h/9uje/kpeHM+0SRS6gGsxnbfmjN6fsU5IdMIP9DcWzVZbxp7mBaaYB9ggZrhlOu
sHp3t9Ndz8kG+ASiJH0DvxeslTKke6h9V3NnF44Ad4kOpFXdYb3YW3u0AEczGR21
LupFSh84XPsCotOroZfmlTe1oBgjFBZocbeVbZzdUjeadMzzSMHtv5VyhXL3sGTN
A1GKzvuNuzbZZDn6Bko8MB968fT+3QCfz0oIaIT7WstSb1y92uZVV5K4RtJ50Hf6
LpmptfIStkMALJXJYvwaLFRn/TEvvy8NqlqpqslvfEP6TzFkGMQNNbMtx2sydH34
XW2m6DWCqFrBH5LYWfp2tLGOZoE1xrZTzh3Mq9rueGAUn+pJje3d1FG1wNXrtgoS
XQBpUFs+ASXYKppeti091kWEJ1CDBI9sbbcsfGWYEzukK7PLRhx44DeI6h6oyUfc
whZLQhOsq+VlJYdWDIdYs5xXYGpeUAc+rUc7LrY5f2CqGqCrUJd3lNBEleeJ2Nk/
VIIwQodQroDFJ0KKowhRYBXDENISsjMjEqk7xziMRhScbD3SZVvguuFTfm485W4D
ZTqJHUcDTz7ZybCmE6cLokOj22+emaakTDXlg18YOwENVZWCrKh1/J54+gL5O8mz
1dF3tqrF55TO/P3y9lgstx0vUKOG00tT4Fdy3FG58IpYtwY2h8TF8PlC+JeMZA95
i1KX11iCB3Uv9+joQ1syl4B1HyhOsR6fvMCTExZDxqug6EicgRq5hlVRHqXu27O4
mc4S7xeclHYbMbYzOPYP3rqcG2dQ2G9TfumlHuTAow2VaUYBCbgwAYzpBGi3Osfs
Quxb4YUzyOJfGquIq3vl+A==
`protect END_PROTECTED
