`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtY2OX7uwrXG8q5WEBrFfhCEsqApNPsvezBBA+eimYpPc2NuUyMIYj7Az2Lk3KAt
LutMMpHx3GeS43hFAch3w575T6LSUxhCLJ4s7cUVvltfguk+ns8G0adwy8DlpJ/L
btePCi8hNxPownpP2ivputdjrR9ShVABQ/zV3KGGoSZG1Hu1LNiIIkjY7t+YvWUJ
1FKeOfvCWLGkjgFPQC2hqOB43jtIfOJUgydrqKlmAG7Y3EYHgQ+Dw7MPXcDhQ6NU
QbsIRPz6co7bHzMkc8RBaJZO+oGao6JwZLVIC7UzwB++K0axCUVMoe0ihxmaAFGt
3ihZBixmz4hsk9DZW0lgqRwUfBAP/e7oPAcWfF/akSiEIAqj3gmKab3H5/6ufpxy
JOA24NKK0XD1xoGcXW6kqMdFdWjYCLzCtSvUYxKcx4GAXIwTyx9G4qoyF8BTp69y
8UEIwxz5Jksb11kyfJUFWdngLma0tQJafZ/S3EKNF4sC3UJKapMXdMxWFb2ERvfa
s30Tv1HplHBvRizO9QvohngmgoqhzuCC4czDjONjTcONRQTxh3LSBLLrdpJRCvKB
zFD55oS+IaJidGGzXhWZdkxvVn7eSscenrBjsP1oySNGcXRcl2svdZhKiRZ0l7PY
Lh+6SWs9a0ycjx+0PvVxNQ==
`protect END_PROTECTED
