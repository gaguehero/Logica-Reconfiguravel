`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwCzzlS5TWkCnSeGEUdhXAscDp4GSvmzYQ8ZZdB9pezyD7OMae6mBv7ErAl3VZKu
KiyA+jr8Y6X/7oePSx1ECgMwCbnr+cbU1JFrWCXYsyvx2yB5Fh3/ZDIIvPNPrI0K
j3D8iVZzRVgwWQEL6tMHvVD+4cxjMqxvPW7LZ3yw9UXZUT/vk1NJc6pIKIRaSkqL
i8qqmmUqFIy/1huiUYsu7wWfevyGZyUN7ZffxxTT1//dAdxCXUfktouVi+mMYI0Y
JP/4VZcuosacks7RjgNAD3FxNkvD8CgAi0RRm+zoLprO39GzT52AU/RRKrzBfUzF
sdpz0tG/s0aFpgK3u3ZrUUDGe1zWRhyAADAo+9IVeotemjXKAwSQ1O+4h9MObE+F
fhbmkGLKMXXYTdGiJZWrYW4sAmSbtBI5XovnHTT62DELpXVKDnABeDvuUtws/ikr
B5b55vFKNMO0oZCgMxweHN5LeWfq+0YyPYFyV76mWRe7p42r2PBPsZXSefkdSmdR
kV7rWbZSurSTXvdvjgnQ95w2BsgU8oUi020kBM8PF7lPhET/QanZnVLTrP2OdPB2
M+pGq0tqXGZ2BGbz8fot21lkoeJKdE4zyiwyHkySWQU1EZuh7fvIj7UhhyuRvRBd
IHJf/G35gYxStmDKv+9igJqiiIMxfq3LcYqux69UYUeH6xC+GDv/hB+xABDaH42Q
H3Ho04rZF4s6iAqrb78XzIJwm7FRO57wuGPfUsxjh/wCO3IO6+QDAA/vS5plDcyO
LCkG65406e36Wcf0984ZvVifZc6FdSoev28PZPytuclq3DazhmeXLFSD0tbYA7uo
Ta6k41F4L2oYdZHKvOOanThP8kHs9fCbx7rkU83GgfDY9FabenUIHdISzf2u0YCD
KVdsPUFQcP8nH7q6u+E155bM4vvoMoP8/4obLnOKR/IXBedRgDvGLrw0Uh9fX7H0
dc5TI4W5YvupiqIma9C7isKHR9xqDM2PtONxzVLc89A6SN0v2oDo1yFmwLbZeSE2
U/y3xbpW0hFaX1CQJZjm245clqlwKbmIQ6cSZg7mGuudWskH2ECpYGDDscL31QxV
vSo3bSEOEodQJacka2ykDMU3+2LcbM9b7F8s/dOYvGk8zDUOV1B4Z+78rIb9QFCg
AVcKYyn8ud+F+8Akyr+ueYOMSpIgTLy5OVLtNY/iJhd5KTYJzDqZum6/xIhSwG1L
VMLDNrP1esGVY2+cvp3HbyjQYKiHYWjkPrJVd2oK/C5tBsNCTfLcng5YZeeXfZ37
bmDXKiTLqoJoaJtetsfVqdd1FV0Xwih9d6dUXzD5xQlqgwFM/5nhIQHPRE/MOeKA
XBCQYp33SqG6tcJEUq3UFej+cF424GgfESpK9xOQQfz3I5MfcxO7ieW0/bvuUiyE
qZOXZoy+fDfsJBSsQFde4ja2vhkn9XT5PMvKR5agEuErGKh1c0aa5ni9b+O5uFrs
HGtQmXpXxSEDOcWXWEbSAwyVkH/7Q9BIaENsrp652qDD1YF/Mp2AAi1tLXXTFe2/
6WFkTpRIBuXnvExnjv1Ly2qmCNUeeUfXyyiB/K0j3br5apTMknboO8tH5nJsqdFs
j+ru0w5Vq7czUV85W+Ki1+cBhlQxjOdc7S9IhTzWsMpypMr5/1eWkjG2W9jy0D30
bYVHYGkk6mOPn5Z6jPFzt7rLMoO+g7OdHdtiKeZ3RcRi7Lb4IDencDb6oCFl5pmr
DCdqSmx+axHdctbqcjg3tPP1FjAwIavccxhE5AsYmkwEaF6oX2/mQfGG5uHR1ae9
sqqHLV8unY/hpPYj7/Lww0fD/D5yPfj6cwnQBTbxm04ab9xam0mZYC/xUS8WccZ5
Fdt9SbMCB2Y8rd0NV/aQ2IuonYgL4q8VT25fZbnu3mSPUCy9S/K+lNAVf7xdcy5a
cQEgPLCnFi8vE1l9adrerAaegt2GlDuDJ8UEQy1/bzpU2lM4l+VlCVIW8uuSgIdj
3h1MWyTPNby91RZrbcbrLxtcgGKwCX09RyjNq1w0OMZhXAPp84Ollh2cY1uUG1tg
JnJBRhvBQiVSSq77a3WhU3ghc5y3+kZDuNfqYtfEEzBvxKHK4H+dDDSHwtSbODrM
/wxaxxFDFaYLIuoY7gmMOiC1JbgQAT8bBdbD+2MVnJyzQib3IBcgwPH8l5dX5Fd6
nCpz1YLjOlCrizzAO/vm2Uq2TcWTcibLlpgUQ1Dfc0cHjZpK8PyPbygEbYQQuEJd
jrSI6+Po2Nte/7DtpDt7MCHeXhKnz9kPR+RTlQaUIxdWR8A6vIitYJqDjVlGzHI1
KkWAynCg1xVeAv5+fvBAzCUhorvo3hUJ9us5nYPajOJGfrPJ9FqQMCds3hSNlJTy
KFBT2rk5X4bnGmfmAdEzS5zoEiwtBkJrHS6BFnX5r9dV9mjtgwgeKnPk9IY7Js6T
8FlQl6b5pZxXBAoS+LKQZ+/ZhEvQVvHN/MiowVVG/k4ecc9dus0B0VsQ2/4d4IZh
3vfTXPXRvOTH3T71vHCrVjQPGCeZ2+HW2vAVnjcKHg4iTvX6D4fs8YXleyHfF4yb
lFXCVuNyUYmBeilsINcitZXwiFLpbnqMGhJEGoMP1anOtokNPS5AXqVXuKOLTbnw
YTWaea7Vyl087aeP/U9NhzLc4/icNBFWPCS7DRXIV6E5hGUI66fo3vud5rd5ioFo
0bTAI7TR6el1URBP6GVnJMvl94W1yqnKKtKz+MQ9YsYDH/5a0p4xro9v6mXqs+uF
LJawJRsPazZ415Imm4Fd4LZCqwi7rades9VUYnidKgolFACGWQbcJRYL113apSIS
DlA/ooBAvenUyo39aR2dsLfeJb9SRWfSPOsEiKFBezTRNyO3eOfzjLBjcUMAX0hH
LR4MxSK3e7JWHr6bwXIYLSDCT9qirjueKFJslJ5pRGETNQqdHuL3lAl1cpJ+Obbr
vMWxNB2XSYuO9p3sDzs0odD5cVNIy2+zvQlSv4QbSm+0aLaqZpPdV3wpM0nAe6Ye
81bc62Q3/nyAA31OkVwGsrCGLq525gt/aI8R/bmOjL2SM9rS9BHT1usU9Rw5y6Cl
dIv5YJRh5Nm+xfRZfX6IzRdqsGhqbVsPgZSSqYXeSSL+GoXNGzYTPxjYVgjQcC21
7NRRtYCOT0iGKggaVoHwYmPWrudNCI/pBalRNQFBT1iTE87Eq59MAvqHG65d2cKL
4y5V8A4W1GrAE05RUtpMcyLLvP7YHnwK5tNRySe827WfDcIOWOGM1H5OBSZNfGgL
K8HHw0hnTmWfZ+MIvjVmkO0ekZxYY5yWWvzp5WN8ojQRp+0qi1uiTBa0ZRA7NJ1m
mpm96CCL7obClZ8pX7CafimUScwdTou6I1Stekex+y8tltxanh4X1bEgRoHeuD4U
nZObb01dW6J2ZM1KqVyCR7WAkbf5qzP2ZpfJYeVjAS/rkBdHQaqXXHk8BN4+S7qi
dCnaESoqsD1uGw0PlBaSGGzV/dTnzmYzzxd2iD7nn3d9tBUFaXbdKTWCy0ynEeK4
Fh6Y0Vgs7wPMLU2TPiT6t5vjKSP3SvavyDVKNQpvPOITYYzKE2NTSOyzXibNOt1E
UIdwwqVwtbahy0Dc4YjXMqd+vhfuvlP+hFtQYtArs5efcx/24zpvkNCaUeqPFCoL
FgiteL1SbmXh9yBTnAvc1QDcsLYOaxQO91eq2F20EttMKps3EgKLynGbWniGMaXs
9Qy6mokkYY05eE6fkS42abzO0kec2abrfM+R0Ej1h/8XjcsEY13G4SlGq5gb5RE4
4AfNCqUI4LlO1nUU+Xu2r5iTFjeylRzKcCYXdRd+qb8EcH0LxoLZTDfYzQN8mwuc
eCYpjODEhGHx0XlM87+zb0q5+D0akfTTh90JFWb9aM40jZAEFPYmuocVLpSNye4i
m3EcMUWE8tmyAorPUoaLqNEGuZtVxYZFXM6HzAL0kmmIGVNx/h2gxfbwng3LtJ3i
GslKOFV29GCb25saCE4nnjsEzdqh+dj8Isx0FV33oIgRA6g0LOs6ouf5p+sbLmDC
VrjRGD4wT6PMMcImnAr/dRxWP9UrZ1dKNWo8LiAdD1nsvAVcJlkMIByNZr8wd4R0
hOF209azh3irlbfRJhLppKR6lkeKHi7mo/mIWb9IJm0pTrzrY0B6+hFkI+pH2QSu
EAR9eYVm/rGJXCpEQooA3fMx3YXxqgYs3H29W1ZCAT25OHBqPSjxgpFsjyR8DHXc
Fd9OTI6gsPGIsBLoEYhJjjH/E/N9yzAP64k9FDxzvQxkA2IdqdZrpz9Mu1Q2k4QU
4wa4XL2qyZQivSNU05mJ0K7BKpcG0NLcMZAENOFEGNqwnylKpg/djgzdUPEqhzsD
YhMpe8tr8wVHGPrEJ+uHojZeXUGxLY1trNIH9fRwzrjCsIeFcpCNl/ZcN+90z1x9
dAVSeGV+nDIKniFq7bEodxrvMUS34NBGhiZYEXeDkltNZmloWyYUyfSnIMIkemud
WiPhn+7BeUN0CqLRqoXkSsCaCz2JLoNqWZjoygL0jKLmEVpoNLm1FNK3RuESwjBu
hcCWvR3NZ235oIqW7ZW270/+3lBGizx+2wUxcsALDpxVpUzXC6c+2qF55tBJsGss
hyD2IyZgpJYBFMN/T4/PW0T005ySPpnOLJd1eSR8AVTyFNNevNUrdDLouFAWYQtC
B5iG9ysPov6Kqrlva/TQOBNCk12vadg2ChmrF898ksVjzBawhSHNrtIy/xk2WxHO
FcDtnXjZUC6rY3M2//id4/kOPOzG6ZCmByREimbzYJ0dU7/6SHREMVqSE4KgZA6L
fyFa6RJssQorQIBrxloRLVSFaVjmpfDL2gGCuL9ShNwZOjvXgufokJDtMGG1fdqZ
8XX+A8wq1cJmaEWoo0K6btlOEhh5Nd0cDFIkyJfgrn1H07t3q7wGd2ufEQoakRII
hjmq7jNI9nEjQSMKPSKxZSwFjQVWQ1PIVtz1l5nqN/m7r9AGGLkoJbALjr2MYE5K
sgCDvBjwrKYdjQuxCi2HYYAMzbdSfe8ncSVLM7RclNX69FqlhjFOTLVUnVoi1A+V
lI/8kKVHtdMe9H4qcHcK3wQhH4mBfkpvnjZJ/BWw8vl9RdoCP/zHTr8TydNkegJj
n1/128yFs5GNS6HYd2lbXUF6y1G3LkjqSpy4gnDKz6yc4/n+a79I8cWb9mgCHd9U
vaDybehNqcqiQJpRgXsu2tDRlg9KVAQV9oHP0uow+QNqVxNrtI3ukW13e5meqFHV
ZwTVtDazr9g3lbX1hrMBSW67AboIdZ0Pz89Mi7fqoR+67mtSyQMnSkXDy0b5GM8W
WbO6fvzto9xHjH4ypyYtcTOMZwNGO3B5ZcElPc7JRCWtCtabiPYvBmYMDEtQEdvG
sq8EY6pg3IVKxsuRX3dMXThSWqf44P8dg2yQpjpQTOXCH2ZI9KyqvXCv/yxHWMiW
9IkUTvB11L87YMsk4dPaj8YHrosi0jef0iFkLRIXOum01MERADjm3YSc8/bkWysI
/f1B0iXT+hs4aOWlN9HFOQ==
`protect END_PROTECTED
