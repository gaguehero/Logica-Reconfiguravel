`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPqY4kb5Lux5csAaUXVmr8jH+y+amy6Ym0IunGdwsZXeF5UbkvJqWB/NOXg4Z23I
/xC2ZzDJUIE753YbTOwi2ghgJqFHKZ4gpSd5vRjQ//21Kxu5jKkM4IGQSIgodBFI
UQrxc6jJA1/VWIWcONzfgBpkTNuRVS4B4rC/hP/n2S3nW3Gf0mzWa/eaJsFi79H7
ayyT11jUg6Jqpas45OiyQgR5bpr7L5C/6eWM13by/0F58xyivO9kM+rxcH9Q6KJ/
tgCjHDBiYcxu8HjMSxTWVZi3OyBe54JUIAQjPCZ2NR84KzCDT/hGrxjxGYs7oFTc
D6QxLW4ogw8H3Nw38fidlrbpXNuc3irEvPPiKb1c/AqXDGEBxAIOw5+NipzG2ibQ
qnO3odtjV+S2hU5UtOy3zWfkcITmr4Ow9nX+YRFgZD1k7E7IosntpJMKDfD7d4ku
+JXASmzzGBGbXLaJtn+xfL7FP/KKAZDr/6TnrmGzgPrB1PiNxi8315HxBXMDdYQQ
dzvucrs2VNuxRKpuRbMWCWiyLVu65fUe5w+WXsGJHQ5lEgVUcSH2IsQhO+kSuf2G
easZySIt8g5cuMnQ8QmhIW5sWAdTu5B9EvvrAShEJwo=
`protect END_PROTECTED
