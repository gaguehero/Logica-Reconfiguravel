`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JFszUCSQwiMYyUu8/MdO7vdM62UPWO00uaDguOhMHxcMz4GsX/tckvrWnByWBav
VYg86JwSbZrRLe7QxNdF7sPt2yw/1itwAlh7NWzITEh8KrmOY4ZeoLNItUBUbKAX
L61fl+zWYyvF2Y98ykzQivdi/4u1frPSV07virpOh8RHZIqRmQkI8aGEsLodI/Bb
xrEnWo3/cdc+oKyh62AeNexckVKbJCCWLE00LkWoZfq9ozAsOwlgOGtfwBawyFL3
TJLQoMgZVcm0sc2AmwbAstGwaM/u+iI8G9xDFQPM2ZxSSUUScjo7n9CDWpYdwYtN
MnFcgrTE7kK3XqN5ed/PZAb1fLXDdY8CXjsHA7/I0pJDfaa18HwyCdv4SjQxgGzB
Cc36y5nglz4nsxgWy9PV0MWL4LZR2ujSdfZJHzrdq01z/AeA7HaDCZz2ndEFOnKT
CrXXRInmCxv90vlwDkpsGSSlfS62DK5Zi7xWNbdsszkxYCBVXqT9XCcseUayMqmh
BUj20Jh5G9HMuJHbT8l3B063IMq5Pk3rVi1ZdyKcItnUmEPnHzfaEo7mwpUmvnoO
SSxePeJYY86GNIPqf4tFI/J0JaEfKv4GRIwB4BkjB+ml7KnlXpxN8YqFmlxPZBx2
mnBz8yNfh4ILalZH7bG1uypbHNGx4+28wsTfiF6iswoF+miHLgQmM+LDbOFqISHw
0v96+GipfwFhREXf4SunKM9+fzuAfvvuDFjHGpqyNv/OlIeGi9IDyToS+uh7qrUz
G63aQiVm2l24yr1/gklLMIpYq699lm5twtameR8OECNAcsNGzx/DFEshSnaJKKRn
dVKBDw1NRs8HwRuel875b5gjqK/rT1yFvdhGiWZnetIC7U8/+YaCD9dHhSayUiX2
lDmhpO0cBdiS+M9IZs/QaYZmyOLIaNjlt/jyQbm9SFJXu/mnh2kLRj5VPxHr7P8m
kY2C/qMzJOa/pBwT0Ggxb7vG6jVtF0bzgt2+AA55Q42lV/1XvFyoQYIqdZjeY3o0
S2wTGbm/gkFGWh3IsTND6xWdBn8PL/YjYc2SwRvuBFscftRm+fjUf8VmO6LyaAp0
Fcp1f8AVRBo/xQ+IlwJOv3+rMUp8NmoXuXqbfEfBsvf96I3I0CNZVjUwH/LI5peZ
1zj9+NoWKTM0yyFJhOobCxa/ECH3JiOZYBlpEcEfJivS0YBwcNR4pxqmhJrlT6el
oCxcBzYxgnspTET24Dm/r7UqwJJGnLB8U1ccWU1MCpqToH3h8uVt/NuqxtcaQdxC
6nHwKq8VRi/zk6RLAw+8lTGeyEmUD4pWXOjCeU1Q75PDxbxL0la1A+Yr4pBej/Sw
YIxRNz/+Hl+pEUCXffoo55R6UIXrhiR8fv/O8JQYP7HG5Hh5mm05wpKp+oqC7739
gfJXHz8Oweu1rmeWrfjdVRhflv9CzoF/pL81gD1mzkk1gBFHcbLe3pw+lespFb6+
+Mn+sGpv9eyLX4xv5wBAWm0s7YaYKmYjJgSSkH7Rf/q4N6b8ojmrIzzsqYnEJCDG
r6txGcLBeSB7c6/lM6Pwjo/hjCTD+0A+EBdG6+kNYdwBLbmrdtUwg2yta8+wcx4N
x4M/74126LcXGOS1Y/goOV+6jcedBfW0fiTlP/q2rBj1Rf/4IprGfycU5a1g+nZP
JSm/YnzA0sGGoHY9VMVuJYuX5GqReBZf6UnrpC+0iLxJJmrDmciqzKLnWl+5ZGtL
GaMF8dmbNXKS6nmTMXTLXMaXe6D1w4nVG5rH4Xc9IYOrq3urrP53QebA6fMGatVM
FQ5blDR/dB2c3ogD0uRlAR+PxXdU/0ZYW4dDz9gu1F7eCpoKr6Mat9Cywq/UCSdR
ytuvjfDQ/B1gAP7NlfQuFDgBZKxWfgz9ibAINRWuMp43h0xs7OkagdWYP83dHQY+
a2oEvja3wi9MYcTE3Nq4vbCrkR12S61dVI9DqJK7PpjKR6VCYEQl/M5EXdmYx+B8
N2YojOmSLbuaKd9j424F/e4xi+XAUSySHKjBO4Fz/xeLfCP1GVNFos8+Nij58ftU
t3U3badBrlnKG3j+D7g2SIAxheA3v31t7riDSkGCh3+HTanl5+GK2oSJe/AINKbN
Pzb8f6AlSSDotgmwIvhXsJSCExgynRJ8HKbac8o2zU16zqysAe41XqyIbvr2eliT
BsVMvIT80BzC0Sy4ZLB/2bPhhnV+3DEoYCU1o1IIxFaSHiJdsb4lQc3LfpBM1fVb
GHKJo4/IMeETwue0+zO9J9Aty3cAukdDZbS9c1QZwct0+vlqFxVhsqn7kGyuuj5I
1p7GM1pF24w+iBQs5QlsDnuXzjQRWArBYaiMl6Vr9NPD7HfrIa+MNluVosAYyGDg
RYeMBMyRAKIE9Uj+Phj58VS8N7TEyajTx7AE3jNzHnPEeuQLhV/F0k4P7yuYz2+n
w6rEarH2Lz8LRZEvi2jNPJMyumopk0ZBkX4NHZWL2ikhQsPAby7kadWayzFpCZM4
5i9mHP0SqbAeco3pkv69KDP8seeO84Fqhn467YzZG5mwviD5rHfr9GkSQLXnNydv
mMqOvX89avG1Xh9zDjjWPRA8VWS7x6jWJOn8scZA1V3mfcte6EkLmGRI2Gg47rvG
VrZf3b+mqXqZkbEgfSiZtRSICdqu2T4JmZnvAjVk4nrb4546ZyQGdUXn05yXdufj
n851U4bVthhS1iKMOukecDX9LosGmbVMxBUKZJhv23Sr9+jCeq2KsPJoXUGo9Ck/
eLhyZtI2MBgjyQxTW/P3/Xadar1WO8hMvytvnn9pp2KVK/Q2vl5ZEPGzXEFPquYX
3TprBSQYlmfDGtKF91ZzrqVxEqyrft5KHZ6gT6ocbeMVkFJVwMlzOY69zI1l2rH1
S1QkyYvucZVVPfR5HFmbLvvvIsf3ND7s9jzMx/K8mmGTYWbw1w4BzIA5r1twtMzX
44tAhlHm5tgsmND3a1fGMWy7mvyAKHI/en4H8U/0xr37x7+lFC1Zt2dfO7Cu+Rdz
ZPyLO4hIT7ahIKSUGtMlJ5z7iX/L6aetpBZACcYhz0H1D5lCAZSAoQpNDLci+iA9
m+wqh83xClyacxKrW+TwxTlBNf1HPN0qnehlyNm0exEhN53RQoUbYZT+Nk7c+4hN
YE1x1fPYOWHYGRj5qeE1/x5fK/mwHHLuByhgAf+j1888mhWpjCWYpbdtDeA1zR+7
13VHT3VWLh5IOmSHfaJ44ZkIoK8YO/cyH8YLjPDyregqAnqCa/pZFWZ9eC80Vtyp
mJw5zVZOAh1MIyMjleT+QnpuDDUBvdFI0cFWJthG6VooPQjy5CvsZgmbM6FajIbJ
h+BZ0G+i90CBSbPEuqcF5p7NMmxRguS7STNo2I0VQ5sgWoagryKnMGHZEL5uEfX3
mS2jSU083BXgLJXzuCCBQsXRd9FfJwS51Qjf8PvddiH/oysIB81X/kLHRUK0EVge
QV0+w2UxKtw7W6hOF2udf0SZuEGwLvE/FtPuWOcoR6BzN45dGI3lGKvk3dWsZz6h
eS7h/LTsNhLmSqeAZh2c6kWjarz3vX4ziL8C1sHSgB7VGRLgmtHRTv+bojGIDbjE
MFSuuTy4wmAe/04erLNg4Dya4dm4bMOg/ativuODETuzRrQGPyhhyZiIupBk6fUu
hZPbesvl+jgtB5C5HggzN0y9m6/vsAFNdC5SR0iIWx/aH4sDZQU2bODEXW6vuY0n
e9Vzspsw/FZXXVMoN8I9QJt6JKwqHjjeL6Vi1VmYeJ7qaC9W0wnQw4wBcaDjz/Bh
CNaciyRQh/23MxGAWySK0afXrf/7Srpkg9UQUlr9kH7qbm84uinwkVXU17U8rqMO
k1v2iuizQY3ah241ZyBrXhn+JIB52ND92AiDxWzRPuHF3T90V9cpvWqXyNU1eIU8
Ab+T0rjlSqkK9Yitj77BELvayl1UjZ3Hg4u2nPnKOebX+RXjQVJCFAgoT0PwlWoC
ZujOoCqvsmMwZF9u0OKGc+VYk3qO7cPqnvcoHCr5xNmxUceE6q5H+oGshZb9o9mg
MHdXar+VvW3nuSTfnQjjBC2QuB6oy3NNR+9r5v/Jqw6z23aHhuRuMabta9ShALDM
6I065fcPquke5UhW1cgq1XlyOGCduVNS1U92uwfQMaYA8p8lXvLUS2Pbbs3IRTXs
q9wmjjiZFSVVRPi4kIRh7NLNyGfdp0JIMA+pnFMJKLvzr1It4rnsZTE78XBcR/I3
cSh9K4rOu+FoiGyKTUZvqHs3kJgHyx7M2WnLEQ8Cpozv4pduv6nQlc7xr6rtZ8xG
wDxoPl13Imma4BVKMVkFU3cFW4JL1/rKH30c9ZR4u8Myb0beRHKMNcLlv/W7s6X9
4qTaZW6XkLRpX9rXiYEwOB4k1ATXkfs08xi6ZrCLdMFL9wp9SXBN/PVmlE9ayefi
uCXauQGI96Svplvvo5rA99FJ9fWqX8vv1yHAG1AkZo7eCL8j0tZKXYSzbJWzgcnJ
sxF7Nqtz05I9xPjdyVvWHW5tNbZ93PXQPgZMbZvbMNYC2eK5JCZfocXEAF30iQR0
iXlXYQhkA7pLttN/q2vAbUGqPfWIqgRiGGVvsRp/exmunUCCCC6xJmEWQ4S9xKK1
laM55W25ZgtufTFyKpiBQvoWnOk9H2Qbb4gKQ5u45OR+89ugIojh9+HYprpINXJK
ptDytloINh6GH/FrWmwjXi6lOQJT7Xe29iBv7YDw8ps+mCYqEREnEy9p865K9a/5
3uQOznSX3THTkZfzqIiYbH5MhRbL5qbcpyGcQv9HNVGGNlQRcIYO1rqFvLLxFJoL
gh1wdEwZWE1eZiEhRg4zBtLaJNJyWhZp9iU/0B3WJB6+mjb0wyAHG+PzQrSZciA4
fga3br4wU03YFT8tvEe6qHzZFAhDyZj5kJRlu0OaKDRQ38URAV7IG5JtUasFRSdf
cmJ8p7mGdyiFSEOgpwA952mEMAdV8dQOh6vKYg8dRVM/QRxa5c9cwTl/Z9Sia1ft
lB+fVTQ1yp1Zd4f5nvcbHcEeP1pSoVvyhjC7XYzmeVStBUECkc2Ha7Niv3CrmhUL
xhSaUjoJk/nSZZ7PLfHU7jPi1mHnd+9ZfsVOqPz0LrbgZ+DlrZSBVz2fVCxtmg6l
cnAQ6RNneryUticdysngwQqBIIMMjmAVrdr4dvlh6fQq/mfnIOYBEYT4JLrWggHd
T0yd+D9h6IUSWeGKtdkWphXmju6Y/GdcF0CaAUoZ173NpVZzT+0ETHsbZpX5soR+
GvJS1gg3LBGTEQxtB3f7YnkAF94npRxh2g+7rSAxsD6YFfSdU4jS4TfXOASgdChK
i7BOfjAW7kCdvTm++3Qllz3MY+0dqn46ZeLWVQFDOHVphpBISjPoyNEXKFlsdBwY
59RH49ogWAdp52SD11l0a7b8C4B29qmTGYJNFEjP8eBY7lO/bgGgjDqckVt8NE8Y
uLP42RfdgJIVCDhM040UbX8UFX/QahCK2Su2/ojmwuxvLta5yUQczubc6p7UkN2J
rLgIS6Y11QmyWyzf1lxgHnTFXWXBR1U3w1q/48en2DPHRCRpvfSKqe2stN/uHWZq
cqi8i+pozMbrT8GyCjdaPky/q64OlxplZQkASDR0RvqwxsJAN/Gee//1vkklTwCg
WL5DxYYTHtpPZmeursycl7kbtpB+/pRvjaafluLAns60bZVeaK70jlo0ofU6EuIe
g2ePOVSRikmjdA6PRSUpidQxmmPraAUYPzo2lF6Br6pizyP/YcnqbnhKys3AmVzy
h17jNu/ki+VTO5hPnv7YgmGr3oVKyqY+MPb5v8hcM9uk8nbP20YGoGt+7Cj5uR3M
ypX4G/t63G3Y1qewXhYa6IB0HweQuxOwRxjE9k9ytbEWdx3toCZyp2Gbi8FTTJtx
vwhkMFS9kP1fIuioDaaR/SHFgbjxOZn/mtkW72czGHpQh1Hft9IFW6Lp972Mfeje
4pTtRoggNq2rx6GCmkpJxApY9BEVi1O/ct0ruNHZYQRpp0kZfAivAaRZKFTLt/Or
nPIGZ75HzaKyJkKjAa0IfsgGiC1ZfzRBeItTV6i83fuMfEUW5iCbsXOvGL1eH1C3
WADYYOik91qYX5bofT5K5Uk9I5sI16BBtlVDUe0vWJ/LMN+c/LBtcz81OnoJ/WXp
PThvoEPi1KJdZ1bu8qseB3iq+HTys1hFEft8PTEZZp6GsjeyOODwRqVHggXpogZO
jI3X0euBnmf+SoaYMYRjGYdrcAvEwW6ZNYRfl6BK4cqaFXl308nMRPW5hNk3oOyn
2qVVYbPwQyIot2QjyDm5BKPTb72QHAaZ4zEfBMoi1/ardEfNBmOH92TZGEMCh3r5
2Pok+lO6b/ceVQZ38iOE7t0E1tLoM+PHKr44RX4DOBWOgV6X30kpBIkjc7XlV7Rw
FyKutCq+0Uo9/w5XoYqgxMDoef94nXqdR4iQRAy2Ah9kla7oNtSbFl+akjVqI1oU
q+e6yEUE5psMPJIisSfG6yb2upFqR9bx68A1FGhiJx/HfNykrTxzEYdBN/C/KnIj
C8lyklBY8WGSDC4qUiBBZHAuqWJosh+W9QPgc5ig7YqojDLmMBj1ZJrN6E2pqPfS
+fOtqjGZigHcEQaNX9MPIZ67wUMttHu/Td82lCnRhuoJEPCgPCqoA5MZQIT0vdY+
Z18ULI7ZRZhH1DvoOBkRxpKbcVt82escTOrc/aLd61M6/ShF9ka1+MRbhHhCn+7c
BjD139nWBT5GgrvBjFVYaalTK9sJnoP5uFnltbNyC9dFX6O9ByhM/MGjdrqpQUGP
XFSh3wd1DPGd3IClaxm9R5ghuP2tt25Kt7alhpUy/OBtbqgqwpIakA17HQgcRlWr
3SayZ5aOOuk1k9cdcsRMOxvKWOCWUbyGYNiiMbgxiVKX3XP0kDrDZOgCST1+9gBm
UwnovsNVg5WhrWbGd9LFX5NtAdYAFGCKGHCgHiclwAl302R4oqQEaAJayhIRqBgj
Qe32SuyZpmlhYX9sBpbZObXHY4r8AdvhisjAy229f/lOmw8aUSkud0lX+y0hOhKP
rtuzXg9YZb5zHFUZ/JPW2Jt/ynw0ONhMlUGfwCyY4eu14TXntvtWCV6r51gPb+HL
fOtTONunfpNQRnxMWVXFRvlWIeyh43GvanVEcAhrppDL8/RDE76vWqSaedi1PDt0
1uqTOrr0E338+EXjQupqk4WUKj/Gk0WExW3+ewnbQdZsJNYK+YuBYnLPY6n5hc5c
RNmQBbYI5fx6/da/JQpXEXfK4uW5Gb9EM7Ias3JwcG3w7xQtp6Jfx1ar0jOh1zli
420pjLi6dC7TrA3cNIYIiIKKeAkyeRT5NQLRhZ3+F+8T7qScaBociPPlTgZYjMhE
5RDWwSEH0Zkjj8hmDimBtWMW2KHeFl39bbhmZvj38f+cWpa3EAYlLdtWWUI1NdGB
8lXTmtJhm/PFB1P8nd5P2U+xeSvUlVkDKiLGdP9S4sjy26kEDYYm7t23QQBLpNaB
mOrUG8FE5+c98tVtjlXTshdvBlVLEr+/o+Np0+Vxr/PWAbwHEXxiNZ/HYlxZfQ6u
BdVmjvtweq2TyfGfoukoZ2nJhIroWrBnTZ+EqEWEvMuFlEIB6Vs4UlCc9V6OYu8V
qU17AUf5OuChBAhSiUUxVbvLXlmLLI7EnfU+ivDGjsa31NEekCVvaptmmnyTvbeR
/DK6bTNGSyszCOFGso3ooUHSdLX0OygceJ6z3TodsO7q8tcy98SPLDPwF6jKsBXA
ywOHWmnauJC6LnEIJy9qbwdeUP+f1XYK4XQ47WpiXUjw84VQjPV6FgNtEZk14jtK
ovnSERRdJFgdJL8JfWuz5ZMU0M1Q+KVVRT4K5ksWQoGKl2aTdpIcwGZxLYsn20rA
LC5d3FYs/zyA+D/NRGsvJblZhLw75NZzCREHJKToCpDrOuvNtu0HWYpk3eLYzxU7
niEorWWA73Uid070nUjRrJx1av6mtgsDV1oQi7Diar/dTcj75lRfAsDHjqTa4u3H
oF9IZsYxsM4hw4RxXdSst3qfW+0Ye2r0qEF4wYag0mmHA0u0eZLsUtWDeqPshIo6
Ygxp6MAIoW0JPcKp8nf8G5nlOTjcozH0qGLD8UBWEhYoOppdcY7+t6pDcP0Zy67f
y4qm8L56vVjyP7iRFY1apnPRm/8Pg5YZ3XP64SusVLYmc8T9Al4U/hgqFtNbhGm2
4B0WNbd+P2v3N1EVzEsQBZ5pLsmFfYwo1qCxs8E2ZT9I+fdw1r+7bhaFhZo4prv7
yueW1lMQIqrKU0MgMpyqU2pPF25VLXIAiea4r9t/tIG/AJKYQtk1BfUxIogBQF+o
gHEGvE8R+0eVAL4QR0mNiUqB9jWKiJM+zZFXgzcg3d/kf5uqWsCBzV3oTYRqEBg9
AGCHI+CqEt1FZLJAXuKL88M5TACxKqzGBL3mtgND35GX735+xbugrQjWPxhTZeEc
/82eHc+qGkPCsE/+/OP/Twmz2+vYurN4Z+VNb1DWm747qGOj8MoLHrLiBZ4lOv+b
ZXE1pvfwxTNEjwTjDITjv+KB8IKAXQlq1PHjUbFJemPpl2VsdoFnTvqQfrmLoJfi
HvRn8EcXbqaMVvSVa+ICpFUUYMVFpsU3hC1SMaFbmiNfuqW8ufyEK6trsjZtn4hH
x9eXHr8OWvAjkRxZjhbeIeioFCG2Z81LSw8fC+f5kXWp1QicM+Op5euQsoNXJg+Y
FrF8QZd7+cvSAbyVfEPmtksFtXJrmgNKj/OLmhWIJxjRTf8p+S0GAxx0SV2zGFWw
Iu31qIeBnUn1GvDrzf3t1LLhZ3PTQPavHaDrDoAwiDy13vfDFvcLIIwOhnsM7S7E
QrRTaLaRTK47wKqueeI3OVSthiUDWxOHLgmz4Cg70kKiG3aH1ztRdXXgTao/FVjP
iqUAlNXBwLvbtgDBstXRBaI6r7e+w3xiE44pB01LNvTp7uAjBmwqSCnblxbj07Ra
0vFWhUY6IJ2SLqpCvhcwI5XwyJHkA0auYSmdLHWMel639AMKc76zd6DIaaJ96nkU
8d98TXTHF+zKGvLigscqPl3f1RIrg0sjjFvIaJDSL85+y/qYDHPrZiU4APXjBXId
dIDiQ0FOCqJGnFtE5FcIyM7/xIQdicRMO5mbiniWzfe+FIOJuFEYgraw12w8ukLx
9uK/iLQ9lId7XAkFMSac3/OzoYXQon7/u/jrdqrY6oSNe60YKsoLmfkYTOkIm2Pt
0BVxrvRi7Kjz/B5eG5liGSHSfLXRvHil6wuPkPHGYB55q4EIVn0eQdXRpLcmzeY8
2Kz2sC/+6i3AZf8oErpk++Li8fUjfKAoLVai7wcuU4zuGC7+XEHZNstn3dPBRz6z
PSVMUHJCOGuP+j+gkusMNpgamo3WQI8K1KstcwRy3bcvnZtscA/7YlCzVuyolrer
n7uJSMT06vzkpjlLpFN0/eexF4DnnbivTlpUBYZwKgl5F3WKYz9w1xwlqfljKq7L
vHyoHquf+GQdQN6+LDbd2Hwnt/j+kdbg5M3JcHi8KLbhv7h9R3JpUUZ0O5TfDIde
s9l0JA73O3hNrNgR2ljb2ZY0NKrubRe+MkR4BeOO4AAoDDtP1sp2enuLv7qW+ShL
VMdk/CPEWLx42OefFq+VQPHKZfWcpvMMxxIKBbfQoLaV5k52B3y9/u2yo1XPObgQ
Qbe4I3I/9OYw1/7wI8RQTltQSwts+euEgSlt8RYZKb19DtqLBR7lTtDDEnRpdXYG
9yA8dvsREmQt9f2XXOa8iujF8SsuKGN3+Edcu5XKlwfeSi+NxHjzbWax7RegVhs5
JDLYs65osoetFEE7TapXuvOgLM11Dcz7eUZt8IAI8Fv57RTGKnlNxm2htl4b4t36
bCmkGjrF8eH8wjlTwl5xCu1BKMoilzLOO72+AVeQaMxbVK5HOsXYG06rdbdTuNKj
adaglDylNDWNL1EWLw0IhHIYEECj3rdJGnks936HE+peP7/ktmddXowmOQNnWGZU
qo5jOdAFWIEbDLlITqC3D0d7ZetCvvfx72qcSH5BMAzgz5+StnYsnD83PcVbscja
juJ+dvKjYbv9uabhLVZ2BrVRXzN2uR68/c1VpguAi70TbN8uPb9PT69vhv3Iq8Rf
B6UlmJQo8KxTREdEkBGqFdAFME0jyAKpyBUJZuyqsvNz6J3k0X9qBfYkQl0mSxVz
K6qfeqztjpZ/PlVgL6b2A/T3yGPvFxporuXCle81w56vpfdOaTMR+Fw9IvBfzhjg
hNUIoD8hwDSP4wGCiOhU6W9bms4PT+DWN/Nji22fmvpZQSc4F7uWZw1yX3iLgcLq
yG8Lw74fOpljpq/AtVnMNlqsZscX/czMjPB4vC0tlwONwIfnF3KetPSwfU6DnMDA
jq75wOR1u8x+pFfx9Cm9m+ymRhsyvt7lewhOMHTMJv2XbeMLk0CQmNgqg6DIVnee
EUFfJFxpPtGc1pFGg+t1nv+pWKoed/dllcDewtPIwYs=
`protect END_PROTECTED
