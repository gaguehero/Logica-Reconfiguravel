`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oGPuFLjcc+HwEJoLdhJzy+3eIAePza760m32Y2nEUZjhE5aex+QvoG0JYQKufLR7
XAMi+K8EXamIzy3BuPtBtLXtsoLtKEwHmXn9ij0joSeT0WHtpcrAKijetAlArIoX
xeNEJAhfQhf2JHSuO7ahwJnx/r813tqpQ15GB8odBfr+v83LmIqeNk+BIJPlrDqp
a/U3Wcke5/ub2U4FOiwdjLhklPJZlSmf4qXCiSeRMbO0deSpu4SViQCI2+HH2VIF
simU720Lhemlj20G3DzivmfCQ+eAKVrP9/FYd3I8ETRAo/mWi/BkIM81OEGbGHbx
W2MnvnoPnjB7OggVgJdGfVEI1Q9CMUjEMKWXRxzUi3Yin+pPtLKb7SeQFipGAW+E
VXhukn5xJvqH+O+Iy8BklZrHNYGO8rpuCx5n6WKfZKUt/llvQNGBjrJXcuC28XRi
kbR3cblIYHpQJrR/d0GaqNOzlYA4ROBGXF5by+6G5rQeEmnPGmD9P180YOm59G0j
XFntjGjKqIW6En4TBGyD9oecX0ywYkixivKNDyrJAy41y8KnUArnpOZQdaF2/EjU
DvPVTj5VcX7HEAmSksBCYPkuU/D/4WnTsOpeaTpYw8g=
`protect END_PROTECTED
