`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6HUb5w9JldLxcKfQcjE0caTdOSDzQoBzAS2y25wNO7LPb+B5M3JPveZt3jsMr5/
Tj0H/mrkEQ8lTjbPpYViSS/Y3PRpZT8QR2kO2jYej4+Pd3raZgen34IPZjRLZSDA
+uHh1RYuasjpSNvAvQh/Vqwp8cctSoFjjn/BLemzoGy1EtqO1cqmllc636rO0dGb
iltRQK21Df3OalDs6AGVzVGrtoF+sBXYHoLsyWMfxTbzESupxkJtfyzej0x8cFm6
yqaKNc4xVV823xX6DZBdyQ2yyAn6aMR+qDVabERDFnzTSIfdfQyxscnFxw2d2kgL
RNrl6Tv2o6281vKjDwRkdkWMxIv0PxqcgAXF+3NM9uNUEJaWhumjwCvW5OOm4OyQ
vc7DA31NyU3K3yYqzPtHIQr1UwRCE6thdcdWUND5D7QS+YpmSo82E/sWTEyNr5om
VfDbKTocleQFEuIhMdr3GR7+Jku6VPvDxI9MuMa7SiW1kto5hIPxp9wcqv11UC3X
ukKb56fksI2Hi2zeaZJa+d57sZsQdXGdS3vtj5Ri9IiZKsNd+IYehqN2AUZicEZh
kA5narTDQkm/yLbEvl8Usbkp4996kjX8QaMzVm531LpJ+JkHwqxUvDmgyhfT2WMG
KMtGkCl3unWXeG8vafQ8ja9G9lk2GFGKKR52K/83QeP8WgJupL+noCiNkia1VaIy
Nczafn/sh5sQK1/qdIFzMsnf39HcZhLqtidBoCHouawAPFHM4kK+w4kCdw2HvUqZ
A24iZSREJ6mi44DNfcW7dkP/EIWuWkK5Zl/RfzqCt/kSmb+zH14+lEeoG724nJXB
CMLzAN9woq0d2G6NLgvIgVsqJ5lqTjvIY1kNXEbCx0IBx/F9D6D2OyJLRibf/AEn
LcZ1ArrkP8ptRnGDjiQggROcGSHBVwMr/2LiEntgCOobNGih2YNYZ88/5OzE0Q0p
VBXbqo3/9ZWvLc3e0vo++71nynqHIx2tMoNjZDxyDNX9icnptlnR4H7O8AGx/Y3G
7mk1nCNgNAIY3HJs6AfHVU9RAT66Pgt5P2ZvpvHAi5MlTsP2WM5xFXtQHdN/jWL8
aCWP+yHTofaZi/SETtITPphedKtnREwm85fGoM6a0+Asti/pP3YDkM2NwWAesu0d
XvoMOViSIdYpXWJw5alxzdcXzezmeVLdnQUEM3yPrvVvC01G9saCmbVtNTu4FG4o
e483p0XxF0voXu02+k0T3iV0W2Cc8oeBl5/WrlEQMeU0qr1noY8FIddLzHM7EHHQ
uOPoE0q1CxK6Z5Y/tylhSlLqPnk1UrG4RgvFHQlqBLUu6iPEfASqNjEtQwYSVupM
5QV0lfBWlDEFaaFqdSG5NG1r3LretOEOr+wyzY/FzUhIggHuupAVUbhjabqhmTzE
NUd415V1Og/UnfibZtd8cu/00LmfRs4M3MEjJTyWHcwBAqxsPGAyk49WE8RiO0h+
pbHvHTn0aB2QnWwLNU6CrGQdWfueAW9vKzoPWTtD/EmzVobBjAPBGjyozCTJTVfn
3YNHX4H4ZtVkaHcY6nqdPTHuFKHWPLe4lJ1XS0E5sC9YpTYaDyWPVoKZxFsMsDY/
NK8FxXRhezKyEQxK/8HWBfRjjAQPeN/IAsx1E3Uuo5dxQXvkYH+AyxmOFWe1+4VA
/83q9AcYuE986z6WR/EBEdy1zLsrQEwQvMAnOQbKRFn7I+saoXvhbSEBiYSyhbXb
MDtM4kCRIWWQCKTXaRD/MeURSA9D82owqokbTxICizwexCs+sXKk3+T4YAtCXYc8
hNtzcWHe1uk3rhA1/Vf5qvpRfHfFxT7JK7PZCfgn3PTU2kmE265cUrhQ+UmNrYHo
LQwbiwsJyjodYL7ZLv3pZPV4KBkb890q+BeHA+/KAaDe9wtyvSO2/lZT4T2y8fou
deYisBYFWKpjlQRC6TRa7s835YCgNhQTHvCM3noTLqwr4waoYO/sVIDEqH1RaWZQ
cNkaI4eE5cztihT5QHo5sA==
`protect END_PROTECTED
