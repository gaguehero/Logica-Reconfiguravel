`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CF4f/0km21pUJH/xdV5dFbsDaDkqqmpP9XmsDyu9jctxzn6NB/3KVmGYeTCraKK
L3BtQgwUMF+m8kU/IHQGjxYsTbHSgaLCY+Vzbit/ZDy5G2HM7xmKcQeZC6clB3X6
785mWcKCyOBhswG1ayfXpBd22dhwaP+VFp/b9QG4WblK56RyQRaT/CD6EvGSV0o1
XtkPDECTJANR7sXaEjDfiQi2tpmi3/xTPp1nm/5SFDcxzlQIa5r3EuD86JjL9G1S
RJy6w12L36xN3S9ZdBAc/3sqmcotvMlr2mFEtblNom4hYtGZfLvxDGZy1yf4/k9Q
8admux7Tb8FkjDthUl+9N76B4OgioURgRXVibnWo34r82cZCOh+atOYYbd4XJEaa
OGfX09JNl5RIoizfEEcc0BSbnvNNeWJx/P1Ve5T3XlCPv+Lz2NTBR5l3iLVzHEph
iItzYB3bhJUnxEZ3DnazApIPPLktWUxhPz20GyVeEABOIsU3Ar4f5qow0HUugi9w
aNQ94C2eB5h/nqVHZGFu7tp3sufEqVpuLsnkv+6I3ARPGdRCu1bOK8UYYrPRJ4fm
0vvowi8kyQVFVyfSpwGngAN9lpbs4YcJYgXiVPQmR1r03b84a7S7TLUxz9fzIgnn
4Iv6oX1rX09kFc+V869tCwQRSAFxdkzvRa9HykaV1b5UpDxM0oPdt3W45m9vcmCv
OLMM4dCIgijJEu09YFptWCD/RP5svokodsvoFsV20dkNZvWvY1eWJX+Rg4h0xC0P
6vEIHU/5qXlS4WTcD0VHkrm8oZce0UIWevRdPRVXS0egMGi+JcAcY61xN9LkwhHi
jFKsBYKW3IMD6n/x2Yx0KI1NUAC2OzsZ1tfFAsR3u6ZDt1/Bvn0XrbLHB4nZN3Sx
3X4Svg0GkIgEOso6kgPmXzrXvgrAiLRTMUSLjbJSnDFHGg+UrFalM4NaXPv3XPZd
ehjgeAV6BAd9nouXMg5IkiMFRm3OpR9Btanwmpofpi3DIT42dmU9xmn9oXVCuOIN
B7JzkqVbnYhtlJZjkvWA3dicYx6bKYqn/Ro82SEdHOrbJethHVXjof730N9QO4Ee
qwrqfKwW0s7DLYOrWZdOVSNe1xP8VniVNLSDCJwhIQbZecIH++NcR5WlKUAvj8fA
0gB/ayiuHsUn3zWaGACX1BhhkTj8AMvo+knF6vasWVM979+FHKb/isoiK5515YC2
kk+DAlHv50qrwPhXATXgaRpk91jvtudO0VELvSXdBjo=
`protect END_PROTECTED
