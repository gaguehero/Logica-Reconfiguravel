`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWrrFEjtLys450U1YKYo12A7+trGoq3dHCCiLgCmbtNzik9fCLWDynkP+aOL8GPX
9W7gGki4PmLnlMtNIOeFgHlsGHgsvWtg7e2D0eXGrshX7mLrFNnfctyx5vg2COzB
S9MPCxr67BBX6PDrnKmw1B07j1wGW/wec1gN6KvzdDH1KDFpDryKyJavzjWrG47e
iMD9CwCMHNsNsrsBXf5bJtKrFEq7dqsAHd6FusfeeN2GUq8qJKQSoyQtq9Fl3KdQ
EbEw5vk47s5pBPWxItne4Xk4R5EaOeF+t+cFA/l55LTjcxk3Sj8SAth2LufbVAni
5XRw/CWy2HwXAaUWdszlA2bL7gYgHFdWCLLe8pk3ITeizM3inff+iYCI8G0vkfqT
kMVd/1zHl33JperkA1iDkp4+aS/pot28tHLW/4dpUkvCZRkgSwWcBxsrTClXu3kk
4eD/PmPYMZblwc3zScfaPYE+zDDe5bUgiKltkBq9D4b/gLWdEltFhWPl+o2Gv3q5
XJqpL/uuTmX1RS1iShrfAns5PIyeEOmo2DBj+QqmBkiF+HmqKeMXBJXA6HJe3M+t
NLYQ2KlaWn921sThJ4/PLymyaA0+H7qkGD1PK3uvEZFitQ8wV6rHkdyDaOdL+oht
NKhRrr7HY0mrGQprTU5rsWx1BM7rDYpVA0Ky4OnCnpvuJGva7OxkxlsQoQaJkb/j
DVbIFw+ITMFMn/dkXuAuwKPCCKMJ/eopIbRzG+V3qvNLTKO2oHvqIN4yKldfcv3f
UaN/TZ7Zb2GsmcDgsNQ2sU0L/mLLhtoWOCAj9oc+1ysuET0R5om8ooHhKqO/Tzbr
YOoC/zv/sajSm/ctFLNwooLWidNXhpms7oJH0T/fkURpZCEERmgyPHV7UHrvtQ62
JSY9tVIaGN8FtckhiLJZWfZNJwYNS9JVxsnZJhVQpO69YlffImEBCO9r0NIJ27AH
qA5rYPbn//2AGk9FfB4ctZCd6QD8LF7H803BSf4ETqHUzHwlMi+FY4prK6+nvDdX
Kacs+vgC7Ene2m02Dz7JjiKUSYbK8PpkfrEki3VsG0KBU9Hk7SIITeuAo1+iSJE7
bDmsx0Ll8oJYyLDX9Bb59k8OqTF/Vu5KMNLfWAr86YkQeiKK73WAUBw2ys/72AUn
sE24mYzSH3lhl3b/Hg0drpM1eS9iKNNKCODQdSYNfU1rNSHRrXEDTYsT4s1cIQQP
KiuEVydJTBykpPlKulaJ9Jn6dOWC+zyHPtHsCBJaa0n3yHM+Z9yFYufjw4YfwkDG
IHY0Kv5x9YWfI531QPT/2SWtRM/bWigKR1zxeofSON243Nq7fK1NbqlktZ/yhfqE
Kr2a2g1sURPIY1n6MgV48Tg2BJOZMPr0I3+CcHknk+AQcdikSUh31TbNoH87pL2e
7eprXxrM5Is6cLCp191nUzyIZrwqYcI+foEMnt2KJNQVgs3+pEUhbEqx3L1hI4g1
yksF9lIstn3LF8sa1vzm6bsaVdEedo0ZMDubHJgQWo/BdE05VAMnEdef4cH1FfPl
8ucexynZATIGMcbTKGKiMp+A7lwPWmXWQ7wxFXrf4jZVbf9jZyPlAgzXTUyH7kwj
p/NtHVdjk32f7mDdMv+OWWeoiI++vJXi23Sdx0MlODJL5PzzQNR1H2oFwTcST79f
XRszDnt4G8S1rT7o8fLL2b45u85yCDWZo5vhPvm1i3qaqTrkq0lJSFst2Jgl1KYj
1YAn/ezD2R5UlGzQuO2+C9F8QjXcTySKHYkfX5/3+MhPoV2Q+u8ErwVFEq9HmERd
kS2UArvS/VndQYW40HnVYF8OebE6UsjRUu1MbkZ8C3CpL3kk9MvtF8jR74yoTwrR
uznM32CcI4sUawJatwUUNx2/Ij20GVK0dgvmLyu9L1k5cEXwCEMqvGf6bOY3I+D0
B98LrN8P3u8uJH2RzCXq9x0/aQKTSxwNlHAuiJi8ID2IaUeDAUSRfr6wsjSEAuJs
21ME+1yAsZwVYqM1n9I9iXK1GCfpr6HzpybBJzT12BtiG7mEcR1VdgfdPy831ebc
BaNadkdreYSYJDiUtWXBRJArfiSj2oL3QXIeDGAywUOrTKijCmVG+X5BeebvHF2M
pTKj19P2XhMAVZGU0BCaVyIAyAMqiIzl7WgpzMY7nxfX5vIDM20GYg9Cp7HSapc4
l/K5xasKsgdiW/9FTUbbKFLdkoFiF5CiUpJuIEJC+kZJEJ8qo3XKO1ua84tKJhDt
0HIWQkJot9JuA1XcOKNRsImLRmhglf0rwjpYH/hlKbl80NLy/ZxWTVb7W+lyqxrq
gc5UHc9cKFWWWZvE2+eGOZ5Wvu3lUb8si3dhi8AkLozQkE4M3zEsuGnngPGsKRmy
GmXTcHM9MFTN/QWPTtHdvcCWhxdu460WSvF+LYbmseRzTjIJV2HnuJ1kE2p7or09
yaWHcpbM4w8O8jUxQ1FJf38rsOlbEWZqSFumKWXEpShaqgywj17vfDJZtwoNE6ch
iE5CDkKeotFLpfWzpDpu4ShUn1PIDriQYcbjMI/ubX8gk3akzWyTRrxFZqOHypU5
rKWmJ3kzwbgjn+mgjfecF8kz1nJn9tRfv628AHX9i+c+5xRTWShI/6xorJAqan6o
TIkcDEP1VMPpUi+qb3f2BDYMVDWk8YdK9ZRpY+a+h5AKq+aopnPowflTW5E3bcwa
u69SC+jEMaeHqB4FqQeM56IqoMkZq7wzG/a1JlYqBlQRpkK+xM4TBVFphZhtP+mK
IPXRaXfG9153QrVI4jvJ0gvyHfPFc3aemQxIGaTrHK5vuD4new2UfWwmwL/J6tVE
DStBWm6zoHOgXhMBGbNgpvnqzkndqZObLhv4v8i1cCDePgtQMQJ67tIN2UAPTwWn
oa6/4Lq3fVoxcDPnoJ5MgRBAMRRuVZWvmpp+8bMyrFZyKxe+IWdWRq5xJqpRohcG
HjzohRqE49g601bgWOvY+LBfLgaTCxDckdbUGKwuwTtSds2G296MNBSOV/bG3oTK
opwisRsdRjAMZRr9q3euKsRMDJ8lnXck/nFHUYJr41mvbAxqKWikhV9gRrN+TQRO
BOf+5Tsh7ud91w2+n5TKP1QDEc7TMDmYJ5bak6H5tDrb0DJ/tIQUQz/HoUjcassO
pwhIkIQwMVQbqYVp8dXqILxCihMwHARwQS7MyY+SZiyA0+tcfcaYCRNAB6vMpVla
bgAMgVI60240ITc/gbmigIgLPOXGlxi1zjZyLJrDWJRCBZ6D0wXYLFpdxtlVhkG4
6X93lloTB6SEVFRKmVhOHqshIuNcsCIAiYdXdbqqyDS0K/6gj0bSUB0Cq7KBlh+C
vGOUuicvqM9NT3ftOEqbyNl/6lyKuDfdI5j6OorEnjWTxE8/cUnyAzo7kR3Ms74i
HL7ljFQz+0A6Sogqf7BwPmFGJmKua1tjbaBMzhAtVrWHHCSNiHTjDbRH5Bqcl1K8
T4nb8jrUm4kW0BvmE+b68ls6W5c+zQOwVLDJzc55LfAeZsB9BBm7kbDIlX/bVpzS
Jlf3ymwYsvzw0eHGuAREMAhpCS/UHh2VKRAu/6FtdX6AlK5HcL7mawUNytsW2shx
uAYnEUuKVJy25NYbjKqOdJ6vZV+N5iZtj/vD0sll7Z5+YxKct8crv5vmeueTe324
mTztfGPMUXmwTRvdavyvOgl88gstRhdyuN9nXoAFQU1laJXCF3cIhHAt9mRLu1Zq
wql+DqiKi8ylTue29P11dKhww0QuDTwslJTxWLEvi7NahN+7ieImsloarGnzoc87
YbW8/rVKoQaZUixpuf73E4DPMoiFl5TrtVcy/jsjTl7c7TenBqkTS2lPH57h0ujK
cvbFdf/igb09Qs+2PxNlTDzj10rkG50rpM7AAV9xksiARMDwxibrV2dI9Mjg93et
RTYcfgi1tt12voCnPuEz+HLO2mx1JJKnQjb5uYus/eM/rzqWtmMkfn5yuT1mKw+u
IWOs29mtFSlxIU+jIxRJGjqFOb7tPw2Ipw3InuFvBXuLdtZYtNna5D5s3Mx0cPKn
qDzE69nfjW9bADvwlKRK3I8FP/o7QpKSscfXXHXPEVOzwmpYG+6iTQb1bXtLqcDC
Qzx13AG5JLQjwmakk0CgZcdQoC8MlsXpAxMq5aSfNkA1j7k7UMO5uaE4176OIs2/
vee+3/r4sbdJQUq8lZAZSXlzZiKkM6Np1q/jhz2DWD+d9qBpJobNHoJBJog6GBzt
+wcU4Y+pfmeg5ozL42uEMGNMW/hPdu2ekuF8sNIAIPEGwwz258lauR2XoduCWfRt
3L/fQQ+pqSGOMVtEeqCzJzlMCzcr0h3hzPOtMJlcEaQxDaAgygrPiRkEE5QgNazC
PneEDo4YpffElskaJq28sRQCUwx0+cJsZJIjszW1Pj+ydsTht3Ga9Fm0uQSUyyrg
uJZhVaKdKeqOZw0PJDw+GDkZmh7vSsCBAuianSLwEXJFQgYb+cBNoopCWUGqQrNk
tbfTm4aeGXYn1ISsLm++0jqUppZilWe6KQtcaPLobLx2CIicllLohTDyF/qzRoc/
482EEbROQy88j+dYmyYjtFBqdHD7Zv4ADBd2ymf+866Wy+E8Z1N9xrsY4Drae4ez
JTxP0DSGKGoWNsvuwo6iKBZdnkaaPcz4mj9+vwP0ULf1qmumMTYRdWtanR2RIKzV
QhrycV4SraLYujWDNMlP4WSkXwKdJ1XfK4BTmr7KmMOi440GPIimfQrM242Qn6Hk
t+i2lFF6kFegk8nqr+t5FWLaFhdH2/Ns+LlDHs+6/DRhQC95OSgxi5KHHfyEAkES
mCsi6VAgphx45M9KvW91RIt4AUoiNC81F2bfvJo0ab1CIVjeiXdcWtEBNuDGVsQ2
5dJxgyi3snV+80CGIhTU02O024x0sgx4DnF9jpQebmMNLGcM/urK0Mrr155vr4f/
CuKIGLScxJIo8zJZ3GvvmWKy7+nJ6OMvrff6ucQxFZhu8U2mOY1RVcU5rWRNl5/a
+yOa/545tVcxipRWidJ24Bj5U+DsVAlIY2T3vJWQs56LG6Bq5+PDm1BZq3RT5jUN
qnXhDOkxcmBcyNHLa9cmgVxhevu87bmzy3j3vULntPlu+fy6og4/gSa0ntzKvqCs
8VHjghaiji4CkQzyVo9DtjRGeUwLRgrx6ryxlm+vPn1O+tEBzQ+qSKsqDEZs0J1N
4q7i9d+U7D0UyKeUdOyuOwA6VyVWcgJrI3Gqeguxee+CVG7zs3D7Lg5xWois/K89
/ZaAJLk2+qwyhM0NXBchPXOSbrqLTtrbveSMoNeKiM06S9lrq2c4lkkqgVy9gEcO
/yYX1ZIA/9oLElGfa+sLGdFTqnx+1NJkO1tx7kbs9TaaK+gRufEdgs3mvLwLR53m
YJ+u+4BZ+h8SVmkjctw6OormQcH1ppmBXiMes3IJL7WPegbt1ieHM6gJRh2ojUCF
g0UHOcF4iTHo70smGlvUxEbpLSrVVRqZbnXvO3o2ayafztQc4cWRiXZ3npOifnZE
+2Q28/LtTWumNiIC8JPJC2L37RpgAPO6MsYdTSwzzxBe1pNe/di0vPY2D+YM5S0j
mj11sN0V7ZQ/YR9MjAI2iMwSqimFQC2tT36lxvsaEG12EiMP9vuQLXXBpDd++bfj
6a8aycc75DDjfr3rkDFjK95vxMwwMAE8xt2vQrUyvw+znLBLLtkQ6kQHNCqmbiJn
J50hWuOqjg0h09dJHiOoh2womC5M4hIv3hg0g3yi3GI/uqiPJAYDoZfRcFLTG4oU
ZZevwJ3YChwHqLi0s7Kz/jdXeFFISgTgAwn/4/+mcUtN0OuZr1KXI4nGspLPMSZM
oMa0l/4MfGpYx6Vns1LCuWoxMg5JYolIZn5U6wBYny2Rh2Y+4lQ9e2XAladrWdNh
Z+x7NAi8uVAGgYfE8m6eOH/TTDF2LM+JgWLM7ieBGNDk2SwYWpwyO9dmKWs4kOGV
k2V+C+pw/gB985wk6ccWBuusQ5QZw2uRZLOUYUNGCbI6UmEWlHb4g8ZeyeSwMuQU
6fIeepXcz5kCzfb+/roCe7cWLRafjcF+vuZqlMg5kSOdTxFpBVrM5aFe4FlJy/Cd
OHIg144HURCdByLChO1ZQ7gIHFlYUNJldWtq1gf3JsZF3hjNWhHQSdNXQZOZ+0zn
AnMzxghfRG178xeOtZMps+9hVTf6bAfgkhkDtanqr6Wlt7GWZcXFLRGKw/iq69Dd
nuRPKZCTZjnP4BOuM/TzToyrkpQzdfLo4+0O/XeePiiDJkrUckK3JXOrkdQGnym4
ECySgqWl7mwnZENk0vxVRgWf84m58TZ4VgApdyE4/+mEKDgi/A44hU1TDnlEjhGz
CLWf312Q9bzn3lb0zv6W079aZwdQPa/NiEF+qk4wsgw/fhGPRu599cUkzIgEI/02
9ss8+TNE9yaK86SrjOMiIyOpT2nYO7Y5UEw5zLvaGERBAwqstkjoPh8ranSRl/y9
fI5ZUxmA4wt99dzwZJF8rDQawtdkNJUwBtEvG0J6lzjrpmQhdJUykA/snlh2RHGj
Tj0BB8lUkImSRrbF4rnalkTeUi3qwfiW4yEV3ZIpaCGxs+T+lvpgxAZc0QcResFZ
LulHySbDrNuPhzDPQQPFKkHexKpsu5VxbXaiGsNZDo25xtvcrvyrIG5XWKCtULuw
l/XTZAabNtxDcZDCpqWK8JX3W1NRJCDNGTumdTAeL6FNb4yasfbeyFMHtAJcAUsG
Z7VAY2/E5+I/vy2mFuBEBmLyvIu2iFYgFwSEmkWifInmpMNx/MeTC5XNL2MrTYjj
CniLQY9AKDqn9JAsLy/FGKgpusNpukWSdOrA6gLg5h/+VwcJ/57ywtsL7FsdoJxH
kwAtrAlrARZ2X8+7CACD/stGxQiKmFrtrBMa+ohMmzbN9DPKPH92r9ahlaLn5Wqh
8xvXZighkTgKBmgkJZEdnBqC/qF0gWjCL7alxHxQWTlYlV5QJDDNOkbZTexcy/dK
eDPQ/Lt2U155aP3lG/zy0AVF4LJOzCaYtJWkUKSWYNUwb0wE7yCHs3naGp/UZ3u7
b13BAikXLDdvS/8KWGqs7xanCS6gZ0LhP2MXtV5/ecSiLd4rtXpN1tso6TvTVzqV
cTYB0EqochWq2mry7AucdLKpRg9aB4Fm7aFsU1f4o9bUTqhx54rcggWqk6/A9OMV
/3H7qDllZInR4/4+7NsFnQKqC2ffmI1RasdeV2zSF7Noj6lQL9xrTzanF1TYUCwx
Thr0Qrux8q7GYc+2E9l1vHCij2MN3L65eJYIxnSMxMft3qkQ718VHGKUJQp5+aHG
Z8athVIp7TyaCUnO0m02q6AgjDFJlLa6Qy0M6Abm+m8vAuH8vc8i4UZijG+kBQRU
EqAsfVZpAW7LUW7aHUTLCn5Ehq6VWaRCrqvnuKau23YzDP4PG+4Rxx2V6fa93PBq
J9FCZ62H+5BWACkV7DR7ai9k13CUICArnnRNTtNUu/Ezosaggx1aXnjwQIFZKsW1
hGNaLh9uUhJ7+GgcniROHWvmn02tgVX3ti7NU1e2AeKFr4MGILolBNivjq4T+k/p
w3c4RpNFXE3WPIu0SM9kYlm1/Dhrmf3kFfXytVMjrjno4UfvUSROw//J61JR+t5Z
3eg6VRk8sEGmkVi7T7OzhEMmaPtaYBQjW33IPG+6WauvfJlKMjWYt1Pq4Pd4Ws5M
72nlyjl4YYJlIiq74pxKgXtWgRAbkuwC+Fdm3ZETPLg5fJTs5R2gEfXDFys2txa3
IRmF98T92I142s5uz8IObi7g4foWb202aYWEcnoB1cDNJ9Ec59guTE3dgwb5lsJT
FN8KQFCfrn1FU1gq8oLRjd8ULmEaL4LwNICBgk+V2NEkUMWDN7W9uaPCAB76W3aP
MjiPLg/NSBH24QvL4Jxg0pCweFPYGRWlJo16lyG0C2TF/o/fJKv4eTJVd5rU5r4p
VaKb19tGePHRssRwRNJ/pxpU5X0L7QihcEmPRic8NcU0Filp8/p931yFBEyveNLp
APYh1KfW/pOecbg+sALaU+fRoDgql0/gnwv4ghjUuzVbiep3YimYIauq+j7yTh/Q
TaeRCjoQJLUxihhO0+gazbOuzA6717QsP4TLvamoka3wsPXstiU6DVe34YLssJ6X
VQHJea/Rz45bCU/Ugi+b7KJRN2k5vnHHXznfWizF34thRMq8c1FOBCTuOLi3U/bV
aAHNYW/Mkuhc798fxFMffglPZwMiE+jQs8wckiq2MzZBWZrEEygl3fyd5wzNGx6J
Hye6oSYFRbFeEi4NDZj3G5JLDu3SoEHOrtNnyGLy4X6QYEr6Cn2wwYAz0iMTOI3J
Qd0KZH173G8EZYYs+pEcXBVOcQQmMLF0Wp4r54XOcfx1RR1m6Si0jks7Wh0u0Qij
C3pcx0amPO48A72YNbaaQxJ0G+DHXps/uwbZEJytmwU1pzWqrbL8nHPEGDCXfit4
AKEUDCpXNNoUbZUe2v6Nr6PAqAw8GFeFx9zIskPE9OfBs9zrIPgf6TtrTRQ8LLmj
UimLZXBuwkj2hhZ6TgzHcjM1cd4fPH1tqfiiEw9kDwGG43SrYk6hJWh6d1wZuPBC
Ygb9wAjSNaoIqvbe8SUT0M+tx/Bv/ZddeOQWEsrarj25rmUmz/iQYWSbB49joPJ8
IFdUZuyP73maaFAqAyDVb5hQTAjccOA7dc8cHSSKWPaDu5M4c6mACKNeA5qmj/uH
kTBpe2+hyYmGJZIoH7eDS7e/7hyxsjGtrv/Q/SV2T1U9xSsJvWWMiht92JjewILN
KgggMadq+68PzPtWvIEAaGNMyPgU3/dAUg0A9EmSK3kj8a30nssafC4idhUz4NMz
FObUg5xx8Eb0XsXAfVFqeLbxUs6W+8Gswi5R6hxck6RzQQMYrLlc91S5o5gVuCIM
f7nAS2Jwi4lB9jijN2hRltLaWRQginc73rxW9lwqV/A=
`protect END_PROTECTED
