`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KK/GK6/cEHmD6JEUC1euAzB3C54n88br9oaTzh9+cT0yQEpjolEkP4SJIWapN8UF
W/KlA7fBf/IGcwQsFbbwlwFA9OZAWSpK0C3ovlHsEJpisywbNPYhP4VT3goZKpq9
mE+S3U9m+mY3ZoqSnfM+KPpyKsl8rhEG73OWNYdHfB9Hak9An6kbygouUDT80Y+D
h1CrWl5TuYhve5iekBQsZdKHT6gkQe4XyQiKUpCmRuzoGoVQnig9TKtcGsh1spO8
s8jJcKC+mPw8AmR+7NyZIPgOPxdk5BJGUa/iqPpLJlDgSnLwNmUlc4NesUJRcraf
r9U3gFPHezrNJxgU2s7054BL2hffkhWIb8LUQdENgRdjSR6ddkF/5Dj5JAGjNSRO
JQk/quHTUzDgk6PQ7bIv6RAAT+s7T54vO5fcWJFjKtBO1OW2ZdhNez9n6NGnEvQR
pQev7aHufqyU1pdby5NJAVq0hluQQp4701mWmmEnM3xNWd72qm0cpgaj5sf7Iv1y
zo8VQ+kiRT6B4bk0xOqf7EZBo6uBwZJBcq5R4g0CHtzjvfFppJLB7HNC5paFHM8q
ka4Psc/lKo6ipP3gSdjw+pPfjBvgYKS+SrU427nQ52gojKRSuHTXY9UFVX+WYotL
ILgBxqHUH7HlB8KjRE2uNcoRG0slptEZBgvctcZzeVe/rCtXu3RmsAv+RBz+549L
nURxnyySEPVQLw+3yDwlvZCHWPblJ2hiKfKmX81c9vWU3CCJbLJVP0Pp/hOnP6CX
L0JP3x9aXCGbbDUewXxEPYPlslP2mpVIhN5mnEzA2JdzyeEWuqaMExjopRpc01U8
9EeRPzOtQrEyeHiHMkLV0Q2yDLq7MYRsFa4qpgnfJFU48PQOxnuLL2BNPGlxdWHM
zcCGNGMGHgI27B/AgLRExZErx2lqr95UWmbTUmjougcpA6z5swsNt3Cd8KK74xQM
1XdLtRVVuiCjHrjp5nf+fhEHwgHnB/NXnc9w3tM45HEWX+wzPjy0kOEvVikQhTJC
fvoqrPEyDfWDikYAkwxumB0B54qS4bEoeVAL3eqBmYxYwZSMccA9GQrhkzKmpWxM
O4jvegc8QpX8pEEP30zAB9Vt3gQcqys4GNpaaz25H+uVbMKAPiTOaJqZ5PC3hDVt
xdkYvOuTFnlDhipLc646vMFB5/geERDrSCaXHo5/pqRIwTrQO61fEZkWix3UEeEc
DK95H0gV54CxqJrNwgtqw2xNK7ZPXKRK4D5GvgzZ37C0VeCeoCyL+eePT22eh9pq
ypG9tzHSjGlhlLVagRoNVePrmW9WDtKTYimP/Z2hG9Pct/BRdGcH9XidMvNCk3nv
H8D16yzo2HPKIoaFM9LllbqDwjcQW9/ePMddv+Jb2T8PbjeqUdNlOEW0ngqhqCk5
V+zu9FBL91RkibkLxdnhOfMlYeVTcZpG1ChQy3Kub39ZABcFp7MuB/fzn3FDYEob
LPeW0lglCxrOQy48vWoyvZLKfiye1kjux0eHQkWer0V3L2q/2m122RXHXv1r/oLn
eSXY2gm/v0yiOrK+jH95lgcvkedBCs5eb4sURHt+JTa/SNZHEDt0LmZk3AFaD1sD
PjBHCG7FwSyDvzKuX33ibNm+/C3BufDsr23vpNz8KeTkMsPGXaa53U0ieQXI9Otm
ckzkUYrHaTlzkDTm4QD+2SnXCzvKqgSmVztLS0TE1SW9JMO39DYHSQ8qzdCTqLP3
Om9jYwVSW9ttc/nvUMMTMREbelpmQHoo4EJ8DfTjbHFolvGaK60QTXbUDgpOzxPQ
iV5uVEqYGdOwXCyr+22zpwTbjxIYxfLgLoflN/kyWzd3XxM1cQW/yFMH1FMFQCeT
yPxqaBdc2Glozwba87GCx3032DWbBwcZ8MFOTduXEr9yqLTlPocy0Rxm7jwDjrhO
SxNhB2q4HLvi3Uwx3Les7mkpAt1pF77kDrancG60m6QwpkdOGVIzZbNmfhGoVjCf
Fw7pEUjWAC39oO4+kI+00SgWI5CWs8VPPSDF8N0LjvmsjvsJrNLgUcHMcCU1pMAp
ck0LmzTtWFYhRAz6UGwC4Sil2y8AJRKp8D1CbhofZ33HpkWC57Es1/Qw8D1mKR4j
FIBFIxdtG1Q+QYw1a9sFJC4PPaqpr1a95+mgvzEWaDp0zHFL1YzpkDQ9ebb4SQSX
XKjfd7f+hr1+LecauS9nTJ4GgkpiBf2Oh61+kgPSbJyYd6jSLpqmkb65SHf8z6BF
bldnM/+LqRahjX3OgYldiA==
`protect END_PROTECTED
