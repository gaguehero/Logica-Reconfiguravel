`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hngmOsGfwShEzOWANg5Aob9hfljYtdMZ0482/0VGIgx2KU97+Cs4An3n5tkoWPB9
VM1p1VgQZrPrw73Acz7KzhdbVlwZY843O+1DvIXCwmpfn9PuTynhBPE+SvQdD415
OukEN7oi5T2VOk48DLuzE1Wznrv8LNmhmeNWa+jt/gO55XPow19iGO/ehIBZOwhQ
jQe75lONx0FrTNOkskHZaVWtjZ1KbcDjM76HQYg3cMeQRne0lpdjo62SzLQfzYTm
b8YhNqYXZRXqIrctyot2QKXpAqVrc83bfwRTS09wWbFgX9HAUbqGLPMIHabyqHAE
5lhRV5v5OLBwkIrbMSXFKk9ReqLRNq3UDWaLmRdQTHhrwDA3aZXzBEjYilYz328C
q6PvnGjGgt9ABMR7o6qMSp5h3i6jvdvV8N3f0A1NNhYoqr1GMXR8kMKSpDWd7VdB
mL81fCiXfu6Kzv0isN3FgAcfJ53+2KCMGX/FnK0V9yzxXIL6uZutwyiiV4RnETYh
93M4jMAwFgNxOjeCt9BCgwmk1S/nC4dvprinGSajR1lHOHPL9pipNVhk2WSwrGK7
VSjUTBIaf0f3bYfLG5UJOzXv0N8itqUfLn7GJJaixn4A0iio+ATVRqp6CRCPJJWt
kBoeo2+fApDR8UiUbXyxV6VjkPNR6ojm10PYbqlwxLvoC+HbwoL7MS+GyOSB25et
M7atzuvYd0VgZkR2WZs6o746WIRXUh9P2u+k4ac0XFPt2dP0ZhZ4Y8U7exjWh+TW
aSthvuCdlT181ByDs2Y+enORe8W1euuK+syizaGFIrTIEKUh1GhONBZwcVIIrIpf
WsP3dVtUyiKkWmacoj7Q3+6EPXRt7MDiVJ005+t1ZiyG1vr2MByKAhz2myakuMx3
LN0pH4g9e9hAtU1brMjpzVcTLLC2oXmVFapmr6p8ys7fBb2Tw//FyXS1M6DpYNZW
II6oXPpXZEE+ntwgHZPoKePZRepHY5rLMf9zt0EsM4sEZBxFBtdDp26bi81eUvXr
b162SG6RSf8xOQrNOJX7oeV08f8j2Z6zUCcfA3UMiKIl87NnhvIpV+TTcopjrdNC
uQfLjGfKQyv0xZEaKSBSUA26GbxWcgU30Q0JCHr5j8UArHjDIaNzxAoLiUQbz+37
aQvlKzX0nxrCzvQOBOKvy1yvKa5bpNyB6293EugiG3XcljnBlxkrAzP4pYjsuY/S
NOVoMmKVwkBKn++3nD6XxfXdMUy+Lik+G9EHJ/+40+o=
`protect END_PROTECTED
