`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SlnA+C5CHJKbwUeKO6o5V49JdqwbxlFCKqH5Dml69okbIGnTUCJCEQ4gdkjLP3St
sjMVL7oTTV71bI/eLzqr3yeEwbI0hu+yY+Jnzokj1KTAaGwwl56S7OetcBXPcT1g
AblpnuaLKdYNEiKlYTQxdZjguEzS2oyt0eD+ftXz34WlgffZHavxKGqi+DR9fLYQ
I3JlO/01ztypaGZuXIWOtUFgQZdji9hNRHS5gprNLffaoqpI592DDhscgAAsTUZQ
i4qKzBTGR4Xeqm/Nn3G1bIyThwN00Lx74AXz92Kf6O5k1Z2fH73E3bDuri0b9lVU
ptHTTBvbS84PyM1AY7VElzmIUlHK3JIwfncq9tscmo8iN+M2rYC2B+SgZyPyz5B8
giE8nLOAFukzggBYdD9//QFhdPSNg/dPROPEwzKNxgolm4w7lW+IyQlD01QTYuZs
N0dHDAWDFxfzL/nk1g0YsHoFgvnMX1aN6UJHBTv4Otl7RPxjsKSrbGMVKjcERDhk
sV2K7R7x3SBI+3/WUW252rWMbheeb9PcZoTD6R0GVywxUIqBG56O7/2m339aqJn1
AXc+Kz12JApJ4bARnSS2/ld0TW4h9aOkiCXIm3LLIWOVjcPXKta8C/PxwqiZX10F
rVfHeJ9vRk9WH4WE4Iq9bzPBzrl27lYbYY9dbY5XzLttVhUQKdQ0OasweRt9CHdw
UyutwJxaCFTCEYty9yJ4ckmDvo53nSHaZqYgMjEuXTYofNPDe0SguwJq7gUdTNSy
iJ+jYZOWv3oFU5R9y76wGGERaiyVczb8MVJeFayxEYRk5sGjHbOznq+Y2ZrBb12x
IsRxrVvSLwDV1z84Zyp+iXO52+2EMl5LzVPZj/KYH44tPMM8LqdzV1PxOZFS3A/x
21nITUmtOnxrr4hh3SkhN4STFxvDFDKwm+/d8iRLVDaUTwVmMhv7CRtolDQwQL/q
udoUhT5eI9KTFTE4eWr6cK4scSljNAFgOlXa1PrSeaQKZ9THb1Xf5UVjLE+uE99T
aVBvcwo7ny5ilhDqawTWZYua5n+1bqy21I+Yd2904gcc2xqzWql2bViZ7ffzH9DR
Cib+D6s+gVpvMpXV8A3gM8kdqbky3BimLjyr3kzzIqHOAqmQmB9kJs5zMj+H05a0
uWWfVSpzPhM9fPHk7y9Vbr3XX34Y5CN6aH8NcYODMOBIe2hKmttCUk47H/AJjEMH
jPkp4q7ik7oS2SLGiBB2W1HTxXaVcY7L3DTIvZS4ewDllCu96JCBjXI0rifBsGUD
ve4jo0h/09kLXR/MiEd2rnJFj+NFaq4N/IWDfuB/Do0cfPphW5S94T9IFmG2xiUn
+UyIX3oXpUxlD+8+4WVjUxQr0aO4RWxVLghKmAIrXJuDo0RH4IM2d4gLuZVQuXHQ
gW0tMu8Z7SbZk0zLjd1kQGMnd+G/tX3ZpeMB4qItlqzACuN9acNcGihr7G4Xi59M
durI0V9RF1i4f4opr4NVT4zjisLFOr16AAuFhchCCn13anyUyDO8x/WVNkfRA9iu
HwJmvMUtjPKfomArs/y44u73ldE3IiKepHcYXseesJBXvu3Q+KtmccTUGSpTyjgq
h6L2REdZTeJduiK/mOkbYWpapv0w/4rvMOtCeOjfEhbUUXP6c2d9L20hYN3/ZXoZ
tcOjV4D6kGMMUS+FCvAt8CGutN19VSNPNwrPPMUhKeZx8r5gFyVMRsF30BDj1hEM
MzOzG7DxKNdhksWpDhqGr/SHTNIp3g6KwOcaXVdnZOy8D3okAK0lKgVs4QAvq/mX
XAeWu3Ypw8sOr8hJ15bzqOWvl+zvdlGU6U22PAwZi0TC41jbTrYDKCO80tbSp5Zc
GzCKmCSI6zo4L+gED6+pPrhUM1m7EOgIbk2ldWvNIGqs6ObuTWpEgUq5H6uHViza
s8bpQBa7gMPEtE1xZqr6OIpyqOuxAwAe7PyDXTe2OpG1a74LclaX/PSrdQUTuImd
5yNC/cIDeyEiZhAmP+XC/jyJfwZqzeB/1zPhO89HqtnQHRc4lNaMPn8Nk9xSIbPx
`protect END_PROTECTED
