`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24Fe5c6XZ0hMJbr55oGpjtLEyKt7E1RDUOUxWiCLH5BARcmEOKGKz0npKQBvIsSR
hyzclWbXCsXJWR/2Q5mtJ3a+Du0Run0fl0mWuYLxjpMLKCfT1Hl4+xRWplgMClzX
uCg8PxpwF3J/IC3bYLTZLYzrhBUcOLbK5oB1HdPPdOJfnj81EV1kFD9us22tfugm
YGZOj0JXlwIunuoxaauKypUs8DGzaDufbrhF5zeByukevlYrtboqYsWahz4zQ6DT
RhNPRDxUHB4FUpGDYblxg9MKbpM33ID/FgwkQKGqxgoBo0dfaL/hUIbQ2a6793EL
DGvfxTA0zU7P2FYh+36wzuwWkPWIGDAPd5KjkUhQm6A+jhzw+Ka9tkBuP9Z1OCcm
bj72W45T1WPcblJjUE9Vd2kwx3JcBRMOR49adFm8NJnt5vOIMlKMqT6OnX6iL7Sp
4OGxi+T44jpdQgwnaY9sEv8o6pL5CQOKywMP1ZI9zRq/ifqGpoehJ2G//GJtUnb3
cKQprd9uMTznSZFfFXv5QMKA95zAyf8dNrzQnQBZWFvILXyXO1OLgy9F7cKLCUWk
uleuj8EuL9SAx3rN6vhS+n+cQ2gTUAZOchDodr8p2P/bbWMCKQ52j6+4gJTEo7FC
N+g9yAnrNeZEMligyf9vWnBnYVpi0Kmz3csG1tRy8IRSsFylOzPY1P2ltOCkvQbG
RYwA1A5c90DZmIMmq1zUhf8d7M0/QHo4UUN+lbvC/igiNmGCjabsNfqtQJWfvP1h
oPoKHioL7pHxYiORUnwyFx1KsVIE2n1Mrd9FMHCis7HvqE8wRDmNxjfv1zG8bZc/
QJ8BJzzDJwjxqolPqpOSZ8M1p664vXCQgxvA2YH6olUYy4O8BWwMiFaTG0b1i73W
RPQXyhB2TS2exOzFxsObrkQRJW9wlvuSvXosGJwDcANhvrsSCifFWtb2JaSTac2v
3uSKdA6resocNbjZL0JrrRDMb4/WysEI973VGELw067+b8+aJCH7ndElEtp0v80X
9br3rQX6smjoHWs0WzR/qhQL/ZCbgXUhHWXuhJ9zg9jWkzAjcDjU0os4cIzRNDxe
AKbcWOLvzLpsarYVAmjgpCcIvAdM84K72+QRHu+1MTmAgAqnUVcl1oQBH+yA8mKu
JWOR+Ac3T40tzUpoen92SKm3cOo8F6oVQsILP1KFK9YVO0tN3IK9bi/0RvpPPLz3
nLYFUgeUaAt/Eba0UndWu/4CZTPrAtxSzn2HSF6sDb2dunMC6+CSdM+Fz0BtBqNk
Y+UNg3GRNYLoeuVjH4Pvmif5RkYZ7w9shrRY+O/aMrhqAr/89WaowR6Nk/VDlHyf
8Nt/ECe5uTxMPzspWdIn4OwWrYziln2iNcsndmQ5hUBwEz4AHUMBPREVyC8NBMAh
SFizOZyELzNzMdgW2MiRzmdq618X6Qe8VVjCb6eDZRh15ujv3WrfjPTIU0ph9Bis
zq4R2RhBW5mrr0uI/C3IiRmbx/E7NatuMSnWy97AE61TmAj+90JdyZpYL8DVxiDM
fbcT9HL8ynKV7XTBLtKGaXgmf9lI5cWPDj7aKbHBN/g0X5nbIHUlf+uCOS5Elud6
JpBMnB6MAejU5cMrozgYd8X09p2/ve53B4wqM+fXA6gySuCYY/qlyyoqTvLR9d54
cJniNIZVAdUHC2JbzRmS5SxbV5gSO3JReLF9La0hXy6eGD1diQOS9ft2bqqMFaMh
PjCdUdeGzsCeUq4rDB0dL2VVEq9hPExXymtf9WqhRo0+2zeNk1An7yCBAxXQjYua
N50EPRRv+kTLZKpigrq0ayFCFI71779sLmyExeUssUUhYyCIRwNh+BGbQVRpDHIS
wsFAFNs+7Js1bt+DAIsk6iFLeT9kYzIED1WcAiuSeF61jbQkxuJsiHmf7+lqRwvR
U52WVLU7qX1eWGhLekibqOuq+6qTgq5hEwDZeXfi5sDmuESXPCSc9RoTfqSUBMTy
TnxG5ozpsPj6z3br1neS8PadiwcWzFpwek6WLRMISZ51PHqsoXhRXxsWDEwzI9TI
xLHQk3pJb6LqoETVzza9aR9lD0BqTQJSVy4RNnIhffxksyLxxG5NF9+C0S/JApIZ
eUPcEm4gJjpQOcvKMSK2NC2LE7w7BwcfG4sSidaHXUk51H6X7xxug6m7PmY0e2jp
VXZLywINN8+QV1KGKBaNIv43SlhbuJI0RryKqt1GbYboM+B3+hd90bKZyVBr3siD
aIIeRKTTCK4Jbu4rUzUp1Q==
`protect END_PROTECTED
