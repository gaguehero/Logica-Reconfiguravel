`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WfegfbOMr3rcFk09Z9O2ECp1j9zgAnO3d9sTA8Si2jtQF0j20zy/zZP9x054E5nP
9moqq/NZqTtr3LKQVFXLjwtOfV5S92nZxJ3EZwqKL/UFfYUt4/NjnEv7DBtbBQ/h
4NxkMwkoBdDEZ5pclcFJ/ICVSL6fZ226weNn9uNSMeffg3N63pPhNFmFghUBUJhF
3D7k6prRY442OI6/Xcem57qzA5sDHciWYc/+ZwSvyFIj9pdgbr99jJYv+4Sd8mZ5
3aO3IS9ciktZlRVrI3SfjlU0FaA9HN58WnCFu0aw/ZHBorWiV4GfXwUVohe5c5/h
eJcJ5Azw2dxMQuMBx6JoQDg9xmFb6la7X2rgi5wGsDROtcIA9Jkb7AZVKhJ0DKmq
TPRbYJa9Tgnkqp3zszF+vQ6G7pq3cJpgYjv4Ugbsq4C8+P2WvUl4wCI8HFGusXkS
KCELHxI5uI4ssllNKtOxiv2/CCoQsR0Lk6Pk10czntaUv5e2HDcZkmbZDkPn3XMN
0fL5Q6m3JwzB+UBaeqZC83pT9ugJmWPyAeYZMw3UMmw+ypYUwEAip8rg9pr5l5AN
9fbfmNK39ZP5KyGtCIaUQcfF6dm4dwZ8EdUiUFgffDjy4nY8Wb8xYx7R082m89nx
WhEKUyz/zPE0FUhJGpqiT04odLno3LQGaVdceNJ3Vn1fml7TpHpVLKvFNb2rpxcd
5mOkIIw/wCvDNuol9E8sAppeboAvfpdMyOJ13TWxu0aaNDjdr3eaWUh5Wkn5NP7z
wzbX5fAT1xp2J0VE899eqaqCnjr4iiolAjlotYiVUfKyERBiWy2f6b0gZvSdL8xi
Ayy14uCLVJURzJK+OId+UN8unnrRO4UFY/rNTCoDconLsMqxgpIxlCaVYBAjBblE
dLsDjXHT49vIHzbh6nP6VgIiPcIbTf8/Xj0bKkqiljM+kBjxgDoqRs2KQg7Ra5mJ
s7FXt8npnYky9V+FF82u5vCdlTyi6In41En3ipYC/u0vRDYN9maSTADR24rjSTdo
iDoriK1zRsKqzdFIiSh3GUyYmbs5aU5iUTZD7mus/mNFCUm6yj01vmRBOQaY0HWE
cyA8gJQaqLRMWVkSVR13nAwZqU4XxlpE2uXcUT9iqHseNeZZZLDMfKQ5O6attxmB
PptXdIrlwmZufLmKZad4ZTVQWFF+nPErQP5yVdSoIGMphdlNM9xDdDwGccRkVKHp
TGU9X1Og7NDORIl9gh+APC/l5Dwz4mhYWAtW8JmgChoUDGZMvJ40P1OKKZLDciC1
O0CCJDGK+31kn0HvE9IEqvymtG6/q14Jh1cnQI+ekVcmfFAk88Wk5GfcA2KUdYWN
G2d4bAHjLrU1YTLu3Vx85vdMSIsKK+AkQtB/LDHcUYn5O5wspF6jMmZYRzX95HHP
XAOBMjoUDvo8EQtkp1cdSAL6WiqWxD9OTG5dycgNY9tDw1tGVB/08rpO90w+WnHW
GE/8niSeb76oRNTcdksc2jGOtoFdquOs8jp40h0/z8K9wllZKjUIDXTxMW3MSQSp
t8TgWvMUUqQMRQZLB1btnNr1luNbcOYwt7jnaF5kA+Z3hjyPA87/i9o+qNmrcYCt
Wg+P0lGjB9WyzYCVpyRY14KMbxzZnnn1a4fTvyhy7EFs4CgaIVgxduGXRL3/bZ0c
yOL6452VPpLTDqXDsHFQhno0iXpxk/ZDeYFtgHJFYy4A/drhx6efjdWLdmtX5NzX
erpBbY7I/UevsKuCtd9QyPtrS1BPvbjZP6eNP1ZAm1EnQofFfyvKqZo16p4iUS8b
qPrO4RF3c9ZjGWEc4n2iLA9QKW/NifEc4qpDA2zJ1AKqj3RD067YaiFNpr0xVb0G
hE0ep/P3AqBsdqcXSP/mvUFKYrJ2Za1DelxcvuMvi8fbF48iWgXzXsboro2bVT/7
+1bApcXetAbJBsqapOyaOkGJ8WeHzVXpykNrCPISk6CVf8IHz37Rtx6jtPi6Vt8T
pgiXMbfEB6wWA9MJYpljWORLdYw/+owD0Ca6U6WomwImEMRoZuybJVygPJSxW02S
FqX4Ke5x9xFr/haM839Wt4ZoH7jLZWoj6bzBLJYGbH+SotkHH7fV2J+RDmupN1+m
0m4e9kmXItqz+sAgG6r1s9cLqGoje85gnA0qKAm+Mwmo2Wz2TYrsVEnfTKtFDMY8
eif6GaTRYcNh3zDGMAp5lKYZZtUMCttWfrKPEOcbzZh0wNivcqAqy9HDP+w5CDrK
yoUNFubWX+hy9kM7ZL/r0oUE3WqCggduAmWpBSoq0TYfncmkg23MNVJryedzLJ3L
eHiGcT5xymHzmeVsYmvWadTKbYjgPB/6fU7k8Y3NWHoQgBVwykUixlvaHGTrlg/v
YpMcaBX7M0zcJ0+6lQFlmO8WnMx+f9napSPCxNvLXhQ03zw7ugssChnLS2sX28Y0
Sk6tUO7bQG86Zho8cJB1oWWXfxp3hyvkCWzAR/HSH6ZgVLt01dmiTvDOuPUMnjPy
lG+uzN2lTstP3pm5pdSn79wJ9w3ycUAmMYqxymhV+DhaEZKlgEVf8D4fe+qHXBUn
TOur6I2gPaog0sa4S2NuECOy4tv2K6+VZtvy518OOrJCgL2GDvg4tw4mqi2sEGw5
Jf+TdjghRxzV6apbGpvlywO/w58XCF/L0K9ooTsA4BS+TEwwHlrSya7++uXUFb9s
cbTcjuHQPlyrUpX0ch4EbUEOyh5HxKIJ7cRtrS4NRA8DB+Ci4UKd7EkuxfbFyaD4
dzLyumZgsAH6FC7LCADO/XOBbYlou6GfxONQWVj3AXFSoylmP13EutIJC6foNuSZ
hSZvjCE2TYZupP9GaLYtI5LlIUsZj6bG6kIgatm5bHyo6S1YminlarqnYCMp+ztd
smHw+xuPfLl0CdngggVUgfTlROLPhskC80Oh+N3WEpCyH29nVCmWV/k1ZrTw3K2J
lu1aoOPWyFzy9YBrHMCQnCzaTtgh4SqJrzUF7ja8pKP0Zu4eNmxvf7XuNEf8IyDF
7gKWbTCAo9KnlQf560eIigS/dwBsSJNDSeqeAiHmio3V0NY225gDZAlYHyAs7bUb
pEOLdRAOxM54V3x/oWNnbzOlk4MPmQdZM2kvUtyvQtjcAnbPJIgOPlMoBot0z1ir
yhIummnRaTr516Ybcmna7CATZL1Ge1PUuumm7EV3eALtZlbVV6ne7Vm3+OwedFzq
IXmoKTyAx3tY5T/dDmlFxJjm4bWzSv54BStk6tHP8vFeukClE2ZY8l5iWYfSf5RR
LwQb+R0rC1fwsRcNxs8M+6gN3rso3qHCNxEWhO5KmjR2GLFU7ekKsIcUpdb1p0qW
S6spFpDZfqDvFaehhWq/TCJOqb14ZyBl9a8ZSOvO4LOScBPRmkBz+X+4vbN14WkW
YWcirt2/Gkr8D98q1r40o+QPcEFnEbjdmlzle/SdoU0A5y0gC4UCMGvnrthPbbHf
MnQQYB9un0AA08l/DDt6kAycvi5eOAnh4ObfkNRubPA9PcSX28iI+xH3fRQaS/sB
+mFlX6GL6XPZbSlA4OcM09tfG7zwAqsL1axwRBBN45sKLHQGBYxx2zNJR81GZXNt
DXf3mp6adrb7dQmuzGV2/LhicO9MUaHHpg59HCyIs47yYLCIRwk6vbNI94W7LPKx
yTxYBtrKNMHtmD8SiGKRMfnhv5W0aq7SYbuvs1D1ZuwFnpBYdeao6C3a8b9iB2UY
Yctn5jCJAKWIfQ8rAgoQSzvMtaoLMfGXRpxZ0c5a+CrfxBDxXfdh3J8R7bD66TCJ
+NhzaUsL9RRnPVGp7PEFy8Rh9HmrfGV+OG0OIglXumyDda82bZ58rvBYzx2ymdHf
ajJIgzoLALoQEH0ZkOFrF+iQNBncS0b7yyUJJejUVPGdtGtNk4W7iNrNzwyiKm3k
BtmCdpyG11gyfeH5xpD2Ie8klKMn0xHJ2qsVqWxUC3REMo4aeHogvEh4bDkNLKs2
TSC2GXV76YlRCX1+Rrvp4qezgBHyOcBed8lJlBqtyuDJHdzzmmmJ5C5aaiL4W7gG
aACflVb+P2NseY5quVJBq2i6yg/mDNqCQISnyldz20NQGzFGfY+Nd7aWbzFjeiNx
T/8qK8Y9IwzqoE7D30984FVdq5LRvOlP4ffGHPs747GYIspX4fiLJJgJtrHu2Bwr
6Upoaqy70JGBP2bekA9Ek3EET/sWzlechws3OSyeu2UWyU1MSTWkaq6jc7Ok/PIh
NV4tntDAD/WiPePLE+UQhKqJDjzptlYE3haFzBgroGhgQc6c/0tHvO6If6ZvYc+1
RH1ZDHCmnc6v4Wym28w8x2VHop4hVY5GTMc9eDyOksudbQl5Z9W+7hXwMBnFXFz1
gTpYB2tkJF/VN1qfB4kzh5XpjLWRoSsCdR+xwHmLwkDPRI8CSsfV+CRmm5E/O3eP
aDPL8OwdkoYvJXfKQB8cIPHjfagSrnNik14aLuBf7wCH/58WXZmhO5lfSXSchHbw
e483i67pvgJhcY5t8JEyLeyOrHE+xQ0lmBsB1BF/x1QsbXQb9dJ3DJwH+J4QqlA7
ecqXy/gxdkSdanO8d8wnMgG5Q+OqC8+30Xs3c69MyeMr525V9EySFe+g+nis4g48
Y4XfMoqcwovjWZgv3dZSCO9o56ssLLEN6qq8/2r+0aU+uX+fkhKm37ipsKJR+n01
NgRJZyEwiK8OkMWw1C/DJ9C8SDkNPzwj+l+EPzh2gSV/bzZ4vSk1L3ycxGMyeM5+
Z8lrMkqOexyaWIj+oK+gEuGEFalu2IdS9UH71RFB5WugJUF90/45CvccNDF4CTaA
tg8kL0WOUrzo8gh52Q16Ivmdve3y9p9aiL3Alzdw9QtA9/n5VicT95RDAvW2/ZIB
+FQ+/7fYfj4uu18ShlfpZaTBh4x5xjgfIVSJBTf42rJuvOv+7AgKVtTqE+b8fSPX
ZKYUVJCDAgFyH34/ZlnhMDxjNERUeI0RWYjlaSVrvqrkP87O5Nh8L9Lt6E8lQBgr
Xz91TOEYMN3DFsGrSqSKjh7qbbRnsPsDB7zEmAau/xjngztgljBaTi7mmGaSDJRQ
7v4XmRRF/LxN4o3UmZHuELm9kPYFXNm4MB0PotFZ47PLljKx4bT0Yvp7yokSPLXL
lPiuxtb8uRPydIZ4A5DYu+rILYzJnT6FzYc+gfrFp1H1c8cyOBPs+B0dZj+6kP6q
DcAc7QMA8S62GDU+IUMhYAqtYivjZ+TBcvwFfLvE8fIw/PQZ/Nat+ZP3Tox168Qb
kGQnAgou53b/XiuiFr4p453RadQLJtB7Bd+ri+Cs0ig8wiHffGW959+h/q1h16XG
eMBldVWyTHroCDsao8Z6z+mLXaY3uXTLZ33ETqUQXlpJxoLSthRg5Jp0MHm1+mFm
DjC8uYdgpVZmP+XINtL4GJ5BQYGGtbCa7nc/UBYYSAEiimX7/lC3kfrtmdGzMHzr
CLq0mqau0vT90kUI7IorgZw5R2nXx2hTNwkCVmajIrEwZmhzorZi7gzQgynUMRN7
3mJsiDAaTO2734YYe6dZnw==
`protect END_PROTECTED
