`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vXWZjPSsr0fW6pKQWYzz3dBEbEj1o3cQx1pNQGjPeS2wGPKNGefLEo+VRkX8QHM
S/cQ7FrVH5aAnC+2lRMVTdtqbsego/TuFHaJV5txypdb1I7VVWIRWddGKoV4LMPG
9qlLyMu1wk0KjYWWISKT09d8xvvBme4HYlu7EfcFmDNZLHaz+KeKCVl13JaNcIRR
aqAyD2A1zMXqfc21jkPOePEYLfMZo9bjLQDJLaUNownQrkhdV7dHB0jx16/iq5Zm
sr9r21HiPKuoTzClxo3D1jyfK76CMmAKNWUqwXuDRuM5AzNis1JmjNozSuHbsLzO
DhJleukfJoAEkq1JCEb7r3PNb+4DhHk4hyDAvquTAj2DpkRkNRvkHYnNeBHGlXND
dEML84//B31F88GxZwCw81axABqRTvJtDkwERmra8eNu6Sm4w4cR/qXBOj7LvYCp
jM6/cvrx7p5t8RFUUF2Uu9ISXdNk2k0CqSMTGm6XjqxX+YYt+gFThbROvCPqQRoJ
oTxnYtPPdUszCbQdFVqN9++yeKygJny59FGaPNjqIXFoIzhOaDN+kqwAIK+EXv2H
n2S/s+SP3kvqraB3i5svo5GcJSgW+x5gzGRRKmsy+ZWKkOnnuPUSF6vaiHv2WvM2
EFIOHxc4FLvWv2efAv2C6WB+YHs/1bKqcKbE2ArFTDbsmK1z5tZAUX/aXKZqtka1
HMHTSHWGoLZd2/We1JsnBiuW3Pw23hgZ7vcohNf5yIb20BfuykEqSkvyCLPaTaY1
QLtab9giphee4AfHM4sHnl2z99kUljHc7kStryqTg0bMD84b1NJ6HyOLytZOgLaV
FPwJ01OCZCySzs+rBkNR4sbRhlOAD8fv0sZddg+5jZBW4p6CewlTdkc8FlAYyTew
O417N6auf5SRYbE/IV3dKIjLL4Sm/F1/J1rrLWzW7nsLrjbti+Pz3Mdxm7/eGUcq
rZXPkFc0ui9bw7sIsK9iEPOxCXey6GCx+FsZG7s2SmgNoBigRoR8nFlKko5m5hTS
dDYXVGcKdAHYDXZFrEJfIG3q2lu84yv8kM7XJUgHjoJk2Ty8tmJh0gAbQ8IyAqgw
06DbUU+ifEiJ92tU97HJLHckOoCq+XO23YVfv6rpGvnxD5zNyVtRZwEjJxrHpRtz
+kJzI3aDDqMemRZ8EeyVKn4hiLvjKmIrCXreHp38eKPRtexp8r+K2g30b4RSAXik
l7zfEKrqZhdlsvR/uKKJ2jhHHBURr0lvJrP2PYwBA0p/YGVdJdsBAvYOz0x1KgDs
QmCCLTj+Cev3tvdsLom+pzBh44NOrbXZ/MVXtH0O6Ipal4L9Bw0X9qdxc2i8M61k
zXr4ifN4NzaT68ksqA4oj1sLjBNJzqBcj/N0vlIb1BiI7Jcs1GZgU4ujRA6FkQU7
txzuDnBj7FtvYc6avMLezWSI64t25gzyjf0L9rfuHZ0V34F049EW9twcmeNkYj6V
zMDzguYu9URRbicyuryPALTtGpuYM7JLdk2gJpCvPsby3r85BOK9JM2LRovI7k41
jVkFYxjDHe/tvzfuidMZlBNn8FLw6nhcItEVqEN5DzfBrXXgHiL6Ehipyef6OaJl
qXR8GsUWCVTxtoefIs/oEAYsSmEbo0Tei3Bvd+0f1K4bsXzO6gEERCJ1vBjKJ3vz
j6MSrS29r1bFok5itTbkfOLl2J77ym6GRYKknBxpbST6j2VrTqfKehzd2wc4tlYE
z9ltEbPeuVbjiIKULWJU2GByt6TasClx0zs4eCBdn78wffJSACklQDxm1IZUaQTV
ZAnDVnG9FXO5ZgKFHP4BFtNQuJHeBC9BfFfGkFIECY+RNDRaSSI+azS4RiAbStep
+SqnKRE3+xsdxDfDuVqhullh+pKRIaT8VD3eX1rq9uk4/SdfPYkMycxF8DgIvmzV
tuVCrR0XZ+9VB9595UgHWWnaAJIClllJ2+L/e5AGNJFLq2o8Mpg94F+8mw2p7Z17
Yl9MfBpmeefE913CCNx1zos7C9Uk3xoY24PnS/B2b1YII/YT67WdmdzY0cc+yunA
1t+CWqv3rt4qob+kI2emBJZGg3Ruz+7f5VairxqvbyhC7dsaGdsLNC3wyLuUaQrk
a7bGQKW1g5WZ3szSEJOIgG2tgvEXzwvOvstowZmEvrDYeaL/i4skIFhpPYXfo60A
pN/f1bTARSOU4U+pNq5sNDQ+LA6ztIMrvXsISuLFk9XUuQHNDjV13QObLGzpjBNZ
GOn0ULeZqd8B/UMdMV74y3mAqFEopvfzCJx4hhQtJ2e8EnjVrMQC+tcJ3XAbhMLo
Y3fb2fs9kEjXm05WmzxNZwlh5jkQl97lFeiB4EhmYd/6b0GplJ6OoGMNG2A7nMw9
jIkC27qTo205v3LfNIIUgN0MczrcwK8UzGGFy3z1NQx4HlsYgoxSCvi/HLZbqjR+
jR1ZV7/1o3dNbf+NnEHqibVHfk562tNJ2FRXUsYiIDucaNwykTsyj1BKo0fu+OkQ
mTOwMYXmd71quELlKqjIn/w4QsBsD/hIrIkVKXzD/EnqwUmPcHsNteKmw1cIu17M
SSNNZXSA46w9fz9F47BW9RnRWhTJ1RvhrjjL7go0Ecg6ykfIruZPCooYgZtN8cVN
iSCOmkfoHjYBH+z0Hio/pxBz5qLNFV/vJigmB6zIU6uRm4KULBh1AtEe6juy7hQk
mOIb03lDN4WW+cBb6+/UsSZwvrrEoyH6Kcmq5CpZSw9s6DdqLNmzQS02Y15bNJVF
u0bDWYEjLWZn/QWk+WuH4RdKIehfwTFYJcxdBF63dhH4FPBIpsfN+23/YzhkE51V
rUZm8WcR3MFN1ibkmqV/k3sC2Gy10YZvqFEaNgDUmD9RORbWKIPYOgQhcXRvkp+v
fYxX8ELXT2efh1I6+nblS6eSdwIJUW7PEW0UFA/McT9iwTQ+ezltUKrcP0lpLFdY
IeRI8EWun32+vO5Bl59vqxahLYMxW7HrCHnX8BXNZVkOwtmZgdhKEMlPi0qGQ6O6
hNvqK03OWCvQeijztN0a6mHYW6cFYzvcubHQyUStBsNWyL9b8lnFRv/eFl5/m+VJ
xJ6AMePGk5MnVNbZ1JBkJ+l/AJ1afUBypsLfqK5uDyiqhzRnBDq3YPdPZUBQiGsX
ThcP8juG6svIVU1m4LVwe9qJ9aMUjq+U4qJS3/I+qKkNrkdXJvV9wEHvqBht2eRF
rKWQe6hzXNryjBVFVcrfvg9f6EvhKvdmT57xTemZgvrZeDeNiT24v7bIy0LxxTYG
xUmodxYMRnJVzJg2N7VWNod0JzJ0Uu9CvHpUyfjjjNsKIylwSWyx2+O2bCBcVp5m
iXnxm7KW8Nv69fT/8w6WdyJkQQHOOxFMeHBtx3YdH4Kz6DTI44G5uYaGtV0dSl0U
Gr+dP2iLi+ApmadmBDOaV6tzKkzQ91a6zxCpvxwxgYhMKiYFLQbXQ6Gp3iiqPxxE
i//zYqZrMEfsQyiqxlfCc2USZU6lywf9YOtNZquOxHF6RRDMK9YxiAyS82Bwc43i
AazlTd/9XaGs5ItfRx3JTu7Mn0DWojJ0lcXezOL/kkBYHGPBEi3MZAcAd5virrTK
SaIDf8nmNXJEKTVKd2b7N4wOduT0J2wflD+e+U4huAcpKpFg5+9yfsMgKXiZpJHk
uy52p3vWxH0YjANweFwkpLf3T4h5TlyFR7dEUkmWwrK401qspI9dP+AkxD0B6AWc
7oLsXOaGlLcX55Ys5MxJSnUeriek77ErPG9zvcrgXVnqlob8R8H2sDfKrvkq1FlP
xLOotgYYpBhvP6FluVzEJ6XZiCqE2+Tl7uwq8OFuoc6Twkv4IEwBd93GZfMcBPRy
iodId/0xi6ylmorwMTkQCBF9J6F5Ry6o/qOT8YyHvfQg9bdIgii+y2wILnFlFP34
zVB0yEPCRt9DthLD7ysb7dmCsLVw7eyGDNROXmDPYpXg89mQ0UnfLAVViBcAImS4
A+d8wQKqlp3sHeNjBuS7NUdWEYWykvSVNq01YJepo1bd3OZHw41+T0xskusauPfR
Xgb2hurp7yQ3mSmzirVAinanpYP1kj6hx/1ZjPO3AW8eeyg53vMYz+RyV0H2YsGi
G4knEvL9/H2CCi2wVmDOioBaFb6CKpLnuZ4pCRYRH80EQWeeWO5TSP4TYUbWLuiL
g1W3yckk73k7lE+O/FfjFS8XWfx1MXKbK5XodB1JE7TCLMCvRBkxGNfCDb8hsiIn
3DarbXVBnkbczV/vr6zWW2ZiUhTNhUzh7NNvufn/oNwf//37gzMZwvhb5H5+P3r+
Xowtcns6aoTLvFcLSIr0tTd+3eMNDdetjdOmbTlmLR8CG0i4ss9Z2O3xlp+3HjW8
3d2FkJTdHuJWz2GJ8dypOFfzXZHTR2IBx6g6XPrX+6j+2d79tamw6BCPVHbpqcqG
87qwD1AP8veFP2w9K0/avRy0Irhv8Yvd4IzbmdATHIaDSfMY8OwPDduRgtj3bVza
Lq4GSsT1s/ULel+mapmk9qoxRT5T/e0S/woHjBVg++xww2V6YhbGehPCfMoc/AFl
IngbXkZ9Y6H91mYHul50FEXJH2oqrbcn6gx2flPO2ZXOPRsLYal+IEYQ/2m2Z1tw
GZcO+06i+voUOapgucGx/2qqZhQ/GWy3za9YUJOEWlFE4RLbX3g7ulf0Fki17R7o
6L8Xw2Rw6JsE/Bit87LWbCTjGYZ1V9QNUht5tM5F/hTKaZ2lxXNEPOgA/9uF14jJ
T0oKANzWfIW/ApKYpUm9uYxmcQDysUO657yVgzyBGDF1Di6vSaw4yEMT1XvpB2te
kDJZAKdH8sktORarqcGqDmM58ff7wfWOxEhYT7CDc9QBP1c00U98S7LicXbRFrPp
G9RUhno/YTK5QaD+7S7jXknszr6beAuO3YxbmbLblgaPxVixp1gkkNZ4uXnMH1Bm
iwPCYDilG+n1EwJmqQuZyzYOd8cEHWuqg6vFMbXOyCDY3uYlSN5kH6npgR3lVIxt
L398UO5L59wqi2FvqUfdzFugt1CPC+IE6+Mb3jk+Jp2MP7xMgV17phP2HhSnRe36
vRAs4hB4Ut3nlyJb1AmQZyXyQoYOQhtQxONO8RtOViPoOc7mKWq3je6/1lfyJsT8
G0urcOqwAzNzEPdLjoVL02UrT8P2M5IV/4Wp0THw4rBF1g92PdT4RzO+Iy2rzzSs
my9dQ05+SPUWYuOMdvV2UAbrumyJHFlbgGoSYScWoaw5Dornmd6yS273ScR/KIAA
6zubS7AGhy6zxuNH2luANRXhZ6f5NJQej2lW62JMpvEF9wjDf2ARx67gExdQTR1p
6OBegF3Rf+25k1Jn1/AudDKV8S9xtSI+4+XvdkoAMGiGC/Tdjy8fz0GFkIaNVWzQ
EkCNM+hK4H1jKXJV1dVWO4XOL2OU+/hf98bLR0zhLZTOLCZ2asd6bev59lacdCYo
AB/bqFX+/yzXq52IUQnrbodlOvF0SAV/xTky5BDlMVp1Fb4ocNnBKOWgoRb23cKP
x9jMuI6MCHsDyomBH6h2ec9jkkiXJ/HS8LRYUCntW60GVSJuLPdfMyO6qGJVfovQ
P0c/NrWhAnI/JMHAzqtyGPiDrccOYpLfL0VQXk/aa6H+tUeZrGpFP/6fyOdJYK2d
P2Iba68/SPTeIK2NIo0xylQGSIH7YRMgBt1TWsnVLrHEsF54LjiUZ9ccjPR6f2wq
8UFZjcVqzMabx2CeWVH97PzeNjG0GA7BZHNkqYVTfjDWjCICTPXbaPHgUJppCJUn
RAF1kMgPq5QOr/w8BG1wevmfaj5X1jj60Mpc4a3xZqFEocakRmnKcnTr3C/SLVr4
ijP8lOCUpJ+XekCx4tcdIwCH1srkjq6gd1SOwCuLAfmAjzpTZCEJ++hrmcsrJQ6b
QVRkm+GHztRi28enE9XgdSk1wV7W/BTrlBFoGZ3mXguoISSTj8mBGmLGroqToi+O
1jczqh3YLHEZHIlmH9NIdcpBdfFyIEOM943QqQVJ5OH5vWq/u5XnFU56txz4Sl1k
6sGFKCB7+DY4nGWvVPDTEt/hT9EifJXInzSbAiSRUceq4fK5Lm2xg50NIlls/1td
2Bj+6eT8Nzvh/nUBbEGtequ0ivOSZZpGoiMMdA7uJqev5WLSblcXB//lWgTa2PNB
5XfJen7uXwWgUS4+guPYKdNUOr3bm9I/sHr3/+fYeZxfarR+T0v1qCCl1Gn/TeI9
nufRm02aXaUETeXMMDKs85eXhswPHS1ONwyU/ZtbbC/Rt3Sgti2gTLqlOpsN6dDY
WbMX4CCW2E+ti6ZiPI9zUlRRK8u0C50tKDRji2F4q2/mGW3ATkXKDgqOcFgGbC5C
ZY9obPD/sRFYY7FRR0aQzezDSrv4Qm0tQ41oihN/D5OPylMRntX+XF7sqFNvmKE2
FjFjRI7rCR4Qr/ppaMXsp3UBYqdY2UyaFRNz/n8K1c5Y5Y/ctngxgiZ7tjOHVSmh
OatrPLUW/1wXLv1VOzS48juDXiXrymwGCMseHrT+j81J53hIwbyFZ9uqWGm+ToAj
ZMvMY8tNHSqvLq72/A1FL+ZWncKrxkDBJNO5DP7yB6ULNPYgCdjxrfGZPrzDu1IV
iFmALl3tGjXWpFPxIB6wco7HZ1DTipwuFVWpCrr4Inmdpck+HdFgUMUONGs5Sfxh
Y+DhioglBWojIUDuTR+XHfe/GNqCLN20giQixc80so8=
`protect END_PROTECTED
