`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LeoyuLkxgLIeBJPNLekWzO0ghqxCDBau12cgSKzzvobFFYS5oCaU1QfPE9w40Q8c
mEst/s9I03Bf/aSrxnhEWosX3OJJgzSpBXRIta9AAlYPZ7PZUnWRY33s9aIc/e+u
/IkiBr6L2tA5oVBJVrDcBTVy/hRak4eggpQ/jK2+tVGVd+62mzCaRZOgCLA7zLkZ
jh+PYQaOi2nAPHj9Se/KUbrz/T0oneR2uWKmsWgJ6zls+btU32C8DXebTQEAiBAY
Io1efPwNzWvdln6MLuEVCHw8KAmzcJYwWfskcFfNCyQM9I50f9iP9eJ/riIgvfm8
8upuWrD92KRoQgOPD++9gx6Se39sOnD/6zvnIGSVFyCwtKdxNvOUqagG2bkpDOa0
W2dgycuiRWbVhtUOz30Co5giPjKu9kgeJJw/Aew1nwSSchLdBYGT95oGUrhP8+fF
omUgELkcg4Qjgg42xPe3L/WD4By/DZu35/3KpU+7jD4uzEL/y7q2gIZm4tO52+vY
F6cYxjqrOCtlXX9H6l5u77P5X5hC6ag3QTBi/BYRPKErAvQPWX73JEJeGyXKDGDO
KndcA8EfIUZkKJhbpHRcWA2uDGZba6P4M9PRdNbomhUg0lIjLzmZQycNF7qR7PgC
Wtmbu78iwrPUJ94NBlY3IdtfPwrPUdit5Zsp/K14UcDTG47au36g/9AfaNWENv1m
MFncwcxQ+ooh7hsTzM/R1/auVzQg8saLX/cq1d8h3+ybjDGztD363uSo7KdfRQVi
E0m3/trFe4+m5geUTRl5WaxFei6fMo9MwQPfq9p2ZHhXugFb/ekjDY3MnbkBH++0
uP/cUhptLWb13ZricSEgTON7+ySKHN/jWnXqDNq659aifux/2rBaCI/mCiQE5fnP
zFnF2jTa04a/vJmXAoRVvtaXk64sv5+rOJrL9yEU4+IETZHDqZpLpwj/NlgU/1Lc
sFwCqLv3ahiB+BmZUNnQXzMO8en0k9WWU5ARuyNso7DaCWnN1Hai2kcXlfA6TsVI
1brjOGYW+y58SctRuyJTA26sR53eca9tR4hYpqpXmNp0oAEpe6swfqnK/YOhiSvG
vdPcr4buxh/D9qLTwI8C1xWQ3N0lg0Y7Fjd/SeuQyl1CqUADWtsbG2PKRVvffuS+
4pU6L4sL/ciRl3dv7kr/wvtNrUU029WbOJDyAF3iF7aPxnM3ZwaSKn/ELTu2Ckxp
+oB2MCUdwbpYDIxxYRH9TRhRqQewsdb8SIZCXSl8P+nCqchBbsyGZWyPr5TdX+HT
CNa4Id9vdtU2BXu2Rf/N6oJ2VrbtiNriuginkekTZB/L7l9PgSxeuvawp1Tu9aX0
IEPkC0dX6halF8Txf875oY7CoFyPMNsLmVAFUSSUeku5Yjnjeed/pwe605uCjIxr
w6Z/14kiC8vKZPhWcvN3HvbugcBRt9VnH605cJxXndxfqFYDiOt/6m/Medc33zQC
kni7nrPDtGOVESnIcBw9enwHEFYvIBk9f8fyHE2AIWKCvzUyvFJhcbXuN9QG7k8q
ctlWhVC9MWwoufu4PVKqKddOnDjnlehvMqJUcfFilMdEVj0pfvY4rhQFKNvaNDLj
kbVAHzjSr0THN9pJwIUhvs5q0LICet1rpigskX6Q5F8seV7WPge9IBc+KoV8mEqm
ow/Upc+Sf76POtfwRgmxbqsJSmjQKKzTrbEtcTN7ZzjhQbe2n0x13FJp7nhGYEbY
glOnWYoNKuNZ+VGG5YJDPU3+ZDx/Ytis8PBuoFli8DC+MQgyW7daPuk+Sy57T9Sx
qUITlNyA0gR7sLeL1d6cG2TPbuu3dN6OLMsMgGXcw7ww44MRqCpWtIH9G3a1gsyC
Z65cZnGP7KnUGuaVv1mmRHpb3/SXL/jfjvgPtOr8Wz7NGVKRzHE6f9RKO18hi4fX
fsNcEi+XhCvsJIlD82YZqA9tvIXLqomYED9CxxpjVZ3+rgF1dHwH/U/Iyfr741/y
knm8B8nlN/MGkajKAaxFx3xorViNS71zo3QiTLgW9dqkGeMELyAGoy8b5w5HI9AS
Bo0KYCF1pqNQGuS4ugSgMQ==
`protect END_PROTECTED
