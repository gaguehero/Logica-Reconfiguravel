`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSDbS9MPV6nmz6vEfaiadYNzsP8vMTQF2tdcBI5qYoD7Hn0pSDEZ/XBm5akYntSO
ngwpt69OitUu721l5Y7STpVaOIdVk3Nsy/w8H/c3J2xUnAp9QgSj5aGkUnWgtW+z
OoOCuuzUmDl/o/7zUYLRhnBWWnhHuNVdZ1i+TpBjFtz2/4UTrsLR//5GafPQMKeW
FNPdkAlX52Fu9rLn2DDxV9+km+1aB8JWp7ZMKsJz+eOdh/8y5R+hkSdEEOOk4WE5
W9JG2WPvjuGQAQpb6ePvSH+9ZXPU0f/+VxHuuxp0BxSk6sV+k1i9LRZpWOomT/uq
gwK/sGEgDBbaz0j7hsZAWJsFqvfj11nRpcJ7zFzQxGa9bKiZLx1ADfLwnxs4VZKR
94EAy33DTRJ4xs7uy6nPQkkoFECrdKI51reRXOyZVdUJBNgjHdx5rZx+mpLz2OJJ
nNoziVWNx5KNI9jh16plRdVBjv/8kxrk/QdVD6+4AIb+RErV1XoaWX8UyOTxT5k8
OczttaHvMpDhN6Ljot3b+JCkwSo+5Bfekkwaw2Lf/CqCTOf0aDegvNMWxUdvDmUc
0Gxef6vTa/Hv/yZbB896TMLPk8I4R3N4MQ9iu86H+wtky7pcWX25P2wRuULY0vEE
ZL50mz/8aLdnb7cty3fb/SPMFwJ4oSczeMNvKrSMNdWYbtFatktKlPrl8LKImxtB
g+9cudFV3njEaCHjmOhAXRVEwQSzWJaSDivwO9aQhIZ6JprAoijxZjS4kssQgu6E
ETJzmnbujW25YysKhANLU/jw939kXc9XhSmKqav51BIH5zsg4SFrPz08OLEAVkLb
Ze4Fv2cxeyuVElSMh4goetbXV028qEkr+o9neAxsqm5LMslU2FzDffg61ucMYvyj
vQoeXfC+ooMUsMYiCi72c49/Pe7hKoocJwL2eFjCtY2QxYzxWQ/xH9TUJ3AV5aHD
KEZVUX/leKfwTKsWnXN/FMVtG7blakR9zPaKR2uAvSfkJ8CQBX2y3i+6bGdf36kk
4jnxJ8Jpu+pnywwAbxrAYA0sZNEVZHmSjJ3ZT8vkT4YkZ2OKAiGtLN+bMxrBKDx6
lc44/D1jwc5bNBY7MCp/Zk3G9Vc623BUxtPhECSz9HNrntEU/jTKyTwgpe4sODUU
Sryz+b5opEgZnROxe04tLKVPeX84u0l/ePcHptLovsVRzTnI62svUKzwCyTH11Y/
Qc4DwBQFA1lZp3wj5sFUVYViUtKf1JenWzhYnYZPbQHi4fMKi/mPOWpan7HMrAmg
jlFKJqTjxm7Ku7xP9O6YfHBvjArmua2Y8J8cO/nXl5jPhsQx7jAjPdYGlws0/8wj
hpM89fnd9EbAyHDr6+pOqAl0jDfoNI5CYzLM5odAt5WgE/YDz2bvo/A/24BKWDqS
HP7P59ChjPri2bcQFDMYEw+dny/dwdT875Ydlhzr2XgocBmMhZ6rgSmNscBnxoWV
ZYcamQ93pkO20sSPxQq2QSrgAKJKPWk1n2b/s4McOCnwk0VhF6yefejA4AhHvtec
O2qKf78/NtCQJPCFF8OD3XBzOH11VN8AiQtJmDIusFALgXKkKUOytYSdK4n4dShB
1AcS0VrAAvWGYfQY30pMlPoimaeIDeU088Oh6X/7/BrdtVqkt7hrxXF/rQEKgSPC
69nygnsUJ0a6cbnQeolcj0ltZPwZ+xksSZNmqg6ks5SHvwU8bJUIzLKC3PzYvnjA
4eo4PD2YN7+zwWo4Wd0kDqmRw5P/g6fkREhxvdNh1qLOImLur2bFNVG+kUtjcPRB
XhxljhVQErga1/x4k7lXsKw3690FLXaKYJnE8xLMOjEz6wrJeXrJyMwPAP9F09UN
yX1Nf+a/a3G8sARr5K7nGOgwnX2vIWvLxgBH1LQM5Swl+lthFD2+FvM2Q7I282Y3
ZvgFD7jkLhaWFOVOtoX6WmqCORpoQqM4y2f5nxICHJ/jq868P095uiJ7duj1xUjN
r8mcSmCzNObOpWA8SDSlbgqp0P4nhDFpXI4hKTxzKAA+lw9EgHm5a1KGVUJGzaDZ
9ZPQY3U7KSSx65Lrb+ziEwN0sCajkNaZIpSyk2PUpTN0I9XHvKQpEp6TjaPno1PM
9NsRkdy9rs/NLRXVcqot9S2TbhEqZTU7ZbUt9T/ZchDpiuSpLgL61G4ibZyzTdhx
tnsqbjFr9xmR1pMCyC/hA4kxq/K3F3Vp01momjUt5/q99ymr/kuQQsPSJ2eZlddm
G+J12Mq0mN0rhIZiJsovzA==
`protect END_PROTECTED
