`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+lSziphUCRGpHPAmTccLlzigPEkFjsW7SdXVM10+aexKZPeM+bSgNOfGHem2dRQ
na/wyXkI8zf6aYnQw7hnit0vgPz+Q48M3Y61t5hek9QnXk9cZIXKEzNA+WVdQsg7
g/qhdJhXwpG9AzbrcEqPpSd/jyOE+yHbBMTJgs8nr495Fgnyh+ZOomEEv45+MhKt
igZPXG3g9E4pNpxrYwPjupZzGXA5EvTbf5Gi0JjwNBXzY/F5qQTtcqRfPYGKcUDi
0HFDGck+kxIvIVBpFX4B0+XvBz3FLAvH/LH8DpjuvjyYlREmkmbRrqHtL2U2Uz2P
l2h8g0v1hLZCMaa6mtVYE0DTMDSG9Z7DrgH8o1sIBoeQO92O1b8r4hveXnEV3ZiO
Xt25MzjmKHMNNrqXJD/NdMMDoyrVdx47lIugsBTWmexjExwyAozyA3J+0EPoL7jZ
3usjVULR2s6kApv8hV6hw3U9lfcfOYvbyIcP/Q8yPVQzOyfrT9exzaeRDtLsjN9t
o5RFpHkvXGdnbvAQoO7yqRTd8ftC/IfJ79Bcc5LNzowthHBOC/UB7ctwoH7soeH6
ZRgWX6oYj5b0SxMbrnxjEApJKzoR6X5VclBvTppNdN/u0yEN998mYKBUqa4+PwX+
yF8aIlR1ES28KFj9fPmUfckXBPr0CWStrH3IlIz1PaLoG6SIAehm3dH+XBQee5YH
2kObBD6OasjLy4GTCAaCrfqBgA4PLuuHq3f2c/uJw7ndaLei6r/u1qGeZMs0mMRh
k+FMebLoWhZJWT0pWtM8QOPmSTorsVy4m7gHwKPQHwlEGz8DrqqIph1y5jC5wjtS
omwNRnQDYGjbz2pFtfJwVy/aDlz13sIIo/hfgOpnIeCrn2Uwf1EiTN5ElM6n13R+
x6l0X3aPYbad85LcD0venjjdXuJ47J/+GiD5nMaLE0JCJSKiSLNRFSpgfeQkXX1e
kkG7YnZmwlRQdO8Kn2E4YfUWimfU1W8S/5Ve8h0YR3s2lHf6NcQ6uoZ8UwFLM8Sk
TwaeqGz9UcB7rDFgkbnpahYIqMsCd/By1WwKUqxq538mUH2J9wI5UyB6hSzyk2cu
6G2q9y2k9MiIYw0vZCqaDP4db6Fq2tS0er16lgqN8h37Cq/KR9iGDdVBkBopVXZ7
senFq0ezBh2RO8ebDoxO1aW/mEsZffdvNNBV0HSDEqrUENPGpg8AI0L4tinbBE59
Qs0LgK5ZjNLD0dIoYKrrLPsnJTKLSXmULyj95JYgfZWDJ/AZQFPmHwGZiN3FO5gZ
ppYRzvYyhHkVh4Vewgl/i7tldfTX3NTWraH+BmPqo6l03I9eD/6ZNJuCUIeD0Z3l
gWX4DG/9okBl3HJj7K8ZkBBF6GSyauIQLBXjZp0dQKz4aiTDLXFotrDE+9G/8Hpl
H/52kcBv9uzm8P2fqcuRSgq9HrPpieDWEvkXWInpdkVmqq7h0VS0veDXxqFkHc59
OxQF5srw05dD95Xe9wjSYqKt5AOnvt/UL+BURr0Ah6IHDoRgwTzsldSW4geskGgX
VE0pfx123LBlFQjLvG8kzzLd60PuzEWwiGJrZSMzIsFGUBTb1rip3RU7kpEPCumK
yUzjd3SiBCwyO6bO5PyRK26ccu5o1eUjCCUXDf1bOOL0kOvgdwC0vJYlG0jW2JxB
V9bLFDerVcRMacayyCVKvPGJuGQy9dPbc9oi+rff4eup4/cFjTnsrEttW/J5tIKG
awCzKoM+5VGpX2JwBfd0fTKh0aSfTBBdWEvQA2PUxEAiqxIqOUF+SJ61mtyIUK0n
Bj3o9AKuEOwPNvKCnCcGrFSvYH/xBNZfAiQd5t7B5RYsmvrztUpXgK3iY6jkBsKP
cZGjbR37c10dv1Bsyd7ikJCmDvEi3vLzF15qWc3X4Cr6k6jYuGcV0lQ/c/sitmh4
FMNBNbat4FGwd58XsBYfgXasPj/SqeLogV5ACfGQFWe09t0TEvkdYqjCrqCLmLdG
YvXYH2eWU3awqH9a8d3+kHRAkxpAw5HdpjPVP8Vo0lNIY/ViDYSHuDe07Lfkeg+7
qvnJCHJoSahdTPdssGAnM8uJA+sWHE6DJHQ/R+XPXiRJ19oaar2EjFcE3A0g+5S3
x0aVJdoDEwOLSBrJNGW9CsRvEVCwW03aU9ka1xLjn3lPPYvDiuJTTBkLZmNNU4/t
RM6M6U3r+U5YH5D+pNzFgwDjEpQXHnChFAzJry5T+pik8/H1HsR3DMFuKBJ8bjPF
K4CtOv0YF6ifHphmUNk4EfIXQ6FKt+yvzH6HHDTKiXrhO21gX+ybRL0V6IYGuQaa
2VT9Sh6dRlKuk+4OgP3c8puah6n69v7Wnsgmd3bBrOgpoC6BMHvUlGtUz+NZk0On
8yUaVJ2rbD8fxHSQKoZfxXoUJjQUaX2YkUMXi4I8tjczbxKRTRmu2l5K1qO1eUl6
c0EK07XYandLa0JzH5hvvhDyBAouN1+r6yaSKAzwopHOZqlcta7f4z4Vv/vYRWzB
+l+DE8UpLGnlqFv2HuEUYS31MvdDyWsfH8N+9JhI3oAOmiSHJBdtNrPqZzxDayiH
Mvw5shRXBKXPCmOMBo5yqwn2JitrReTztnIJLPm9M2sikTKefvHoflIeh71IuhjF
eCFYaZ25YhmNAydKCKbEsXVPGXnlumvl1RsEN2iteE9mNdVZnWrZ6THbS73MvIRM
KdNR+1Dme73L+WT6G0fHDf0YI5CNFhMoYcSab8ZeeppTbsiL8kXuM53hBCLhLVVl
TQNoYmaDYxBzE9TiS4fFPD39WOKNnTOHHT+3jAaIkvI9qLGKShtC8veRT/8mepnY
6dRoFWmITnxkXO4oC5QhCRwrxemHbPOylYgXcEPh24ob7mX5bSsp/GxgTGUeF/8q
9BlfISdplHYdX1gKfR6nSRtVYuh39ZOQr3otN3LpBunq0OeGdasc3Gcd4WQU7VAK
W72o9sdfm4KyotDW2UOKskUEpTZI5uDpRThtVidSUoduPAn+6g/V82Zzh51osX3E
oJiFqTMoUc4UCRdOsA8Eozz9jWQGM7ZrQUnIH1k8E7dcF4cU55PqpkiZzeAvrxZw
KAcQMwIZGgUHaaPUqbX37dzF3ESS87cWPOspRWf6NK2TN/HMylGr35/CqB14yrVB
8NxM0q7Z8+8u0sEjCcCFa0me6PrUH8BzsM8vz2VwSCfFPRo0c3tkW+ckMGoIGYYk
dw9PcD48dG0iye85huUiEg/nA7A0/9chYG9ru30o7KU1FytKv4YHzRUglIEC4s9m
QpVRkhGRDYL1fjr7mcJA5OWughBsK1NT41W21wRnwvDNf+29P1D5sGy9KIx/UNZL
8xTnHZoX9MYDm9UtbUz1qrFvg/XTA3GRDY/zaGdfPDlf4PX+l/3ybGc6h+NbVBc2
IemN8MGdKkZW9OmkCTb0iYN46XPh+0dXU+AIDNvuIiaTwN0af9iy1DTJFUDqNxPm
Z3tkMB/YX7aThSs+fhnjQuV6jnXNcUUvg4knBvK+NESaP6lkpLq6HSIPAXjluj9j
ZJP1wyJptp9bB4KmBkT5BgtsZnde4+7VvTMDk4PS+sRVI3Cwlvl997m2DUh0gyM/
W18Vm1MSfisFr+2oQr+aQAhgaFhS97SEhNwiU0u1L365hTphfd39X+sCUWtzXNh4
grEaruCZ3c4gNgWDjcfRUaYpYbLwQgMaFWeft8zQX5d66zSZJ0OuXqPlFaCPi9kX
P5UoVXr8+l4YPRgXZhjji6aohDuPjygJOO8GP2y3BhOlQkxZ0MSBXgsMMf+g9SAx
4qFjzK11oi1sFshDl3S6aj+k4BnUo6JomlBPUlIHXtEoaWefrx3BpDFv+aXBnQgL
DRlj/fziO5GsRObmkhyHDOfvrXmorSNOQUV5DZG9k1Pg5M9f7roNTdQdHCl0ZEt4
DSIT8MLwRfu3QPTqrez+2WaczJXaCUDvvvlw0iTTc5bT+alaMhS0ArLe60nVxIm2
sRyCvJUcfKaquOi0ZlQuchMYyLVQ6z5yOwS80P7H3HprwjcRpAuEcjcRo8N3557r
2Fs5VKihwa259iGGXpVqubQR4QPpf2EraYlZIOSKlQ963qlUj8uVuZRsEpGu9xEn
Fnv62NrxgUlKJQi6pcmwCC4wBuyrm19Ce3QEjG7RlRvjXimeCORtGXBDpep+BhcB
c12bcc+x9eT93g88rYJ56gymtM68yL+vN953u2PF3Cob+J9WB0POlGJ2t1CYuNfn
Ze0VKiqC9lXvycC+kOCilzEpH7R08cTmxVJ2/KGc/rQK67HZ4rHHBBHtr9vV7qZu
KPNeR/wj3nClhMuNbbSUC/U3mfYrY60TGUUqY3875qHcYtev7hSU4X0MwTlMTiYN
y7ab1SVilgy1fRPL6NS31vhKmziyEW0y6HyqAMsK7coRFJZkQylQ32F6h9jUHjzG
QzcTZNtvtjGvD1nb9EzjVD9T4S0ToR5Qz8B2GifLbP9Y/GHQBFkgNrhQuo+VHd0c
nMfIcF5NmfuVEHd45/MNpVG51jEh+OqEH1o4SzHbhCrSdhj8x/yN0xpEAh49Uwo5
hnsg3uIXftulKAHmnf3g/rTeuJIBVO0QnNZ8KmeEIjvnQ2PfxVOPDU7zcLqfUkDw
gSHgTsTkJ77i3uyoGqT0D4/OF1AuI8i5bPWJdm7xbFmmg8ffIpJT4t9QoKfQFqDl
nCjtiBHRLCrNs7ph//4McWnRZFHjMyFujY29ig5yDlnkTQaE3+w0yA+2z/OLk4b1
bFIIbzV8q/ohNN9vUOySYjlMz/m2tCkGMQWHofbB+9P9/tRC0O4VkbyyoWXCzH/y
/E7HJ1KHTZ+q4EQJ7DMu/MmLN+2p80TFSXEHRPBd+km/0Nj7LaV93x0p7bNHDSZr
HHnpFf8Pe5nWDsU/oqNAfYJx1+dMt6XgbZAqJtOo9ezgzpGQzo+ahxkljfyJMRic
HcNwpuSAm8cReHiLzu4CxznN/7foCvFkBNJlpD4dHfX8UV/r3Itygv8WnCXwIMe7
PWNYN7kSIEjVWcSRaM4LiOki3R7FKpjGnUvq19NN+ECx4FBCDqNPQBpC9F0IqXkk
5MYoYeO2gXJydDNlImOQ5dBz4ddtUPZe5gUVwYo+GMirCtLGKuwyZQCMHYHREebf
JAfe+by6nsMLcjkqZBSOjoS2elpmqMe1lrpDxs9NtDQCKDTGK7jWfvfZbMn9/HnS
auqd/ZkfWvITlMjPtIX3cgQE2z1JKcyYKHuYiTzwD1WqXbzRB8C2CkD1YAXpKNPz
fAXljlpueIUX/RruQoiduK2UbPKNeLQ5LSKpc60ZTxfh4t0j3aHLlsxVZrCfY1h8
lod8dMYvC3s0WgYXiFsBuoHseWE12aNU4f4wEsO/3Xqd2A0+vMj8uaxC6R8k83B7
EnVo8fee8vvpBboXqBNg8HgWtjDO2zMUHrKoo+wwXo83V90qJ9FZQLaY0lEitxCY
cDdlprbdQBCBR9kn6FCBd8FxUQteawaCmnCqTkTstZPOBQBE80vtaJ6hPDaJwMcE
IM8msR702jzfTaDx6SsaPQ==
`protect END_PROTECTED
