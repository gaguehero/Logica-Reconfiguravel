`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7XaVwlQv67On0cLlbbDzHzlSpWYvKHOyVGBM1TsFx5r0J5Njv9RWE2rZmBVmwgZ
I20HSetFJeKy3WppvcPSYQVsN4AlwNzb/CQp6SX6USJQ6t2nJImY1hnHta45xGOs
aVv9c6Le64GuHHzV9MuUusTpF9z18Js9LybWUPuY+LOlNlvIha4ZV/BOex4Fl2ER
1R8w4U28BWBWE6s3PXqfK+L8reOlP8BUUkjWrLqk63fdhjUd1zYlVyBUfmOUTfwd
QeCUP2qxUIfb5UiTC8xvFA3r8T6g4PKouBGQY4gTJAzP65oMGjrJIsaBWqDK66ww
l5hJHKQTGBowkLwYUu4zZaXT/g4m+EZf70YgkrV1VQttSwof1v/ahjoSFuXp1bzc
qnxHGqZL69SmR0j4Lh57jUdzubkl7ounW47jPhHvDqQSri0wfppZBPvk/yR6kCGv
t2bqIG8OntMkkOP9AyPJm7/5UJSIbjQs8xvf9w8+N9FswcB2DGMVshqUtK24YaiW
GLawV2s6tG17JkFY+bsb8dWHU1zLYrSryMU1TfjaeMxdXK+6s/OpyW/C8KROnxLr
a9cx8thspS5UvTDfJPic1/IkQKsLBp0kxYZb2znEoj0=
`protect END_PROTECTED
