`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucKDd2oxSxWotbRI7cLYGZ1JKyiPJMbYCd6TjFNKUGHbYmngFtEhPJkfrAOnJfwj
4JsbHchdScoRhrTr38PEcEagcDPzWNfFqEG/lfZG5UtOjHNJQ2erGpBhiLU320c7
32nTTgUaOPw04hLufztdIiAPGYOA2mvi45VFPiLi+IqC8h09ZuzSVWuZlL969tyT
vf/RIiMCAAjDEMBzsbRndhKbm6oMOlZuZ09e+o80cvmqCCZ9DE/O4ZH9PaB30p36
kRrj4aRq8G5m+0BvZh+PzqvdQWbV+owob9j8b2SZ6XfZEqMClEnbb/hcbk5AjrSA
PJUMwPpoutokRgO0FayiusqmDD45V03K9jtCgh3OCIieDZYdIsSKmNnQjuN2GN/+
vQsGybQiD85EmHSG8SPlH2EMCuf3acDEPV8v74EWmAGjq2GLMpjd20ehm7NNfyjg
pe5OFyvM98DC6Rya7r+8f8mdgDvoQ5QO/eIE1lxQinaFJ/tEVstGMtuMpGj9TjQH
Q3QHobI2cqxwy++FqZNkb83UBYWQcspxj5zWfEXlC8G8ZvRyMVRVOhpq8IUrFI5O
XyOYOfz5GV0PeQ5GEFXE0RA4X6LkaVeBYBbzyLtKxGHWFbs9IGj8pH7bVL/PHv4W
U+g+K+8SmgSWoR1jEdP0amx2gHF/4dfToTtdCiWaC/FTOX5842bwTfOJl4FIJEyG
eFUdTDXux5TW8MYvwjnb0GajfWnn79zIYC1kNHL5heAaaHnn5SvF8+KLlpeCxxGB
cOMfG5AZM8AlXjTRqTRD2z68VXTjjMr/EHbJT4dA14YmKwp5KrFpuX5qM2vGa0Uk
Mvgs6e04eDM4T6py3Q7bpQrgcPaq/b117IDPBj576dhNnVifJRqP84sFFNyo1SaG
oKqDwHs/yyfrYBEtkF7v3yPCahaxOb16pFcuEvIHGKhO1o1j3jcrF1Pun0Uc0ORA
LXiEKZxhJ+cAjy7KGXwH3EW2X7taqEz7yVXIupuZd1ykjy49DwpZd+cWgNo6nli4
rCWcnih+qpH2uXoEionEke9Lm0WfhxQFEzZ+ESdby5VHFY3JjDGLGVSZS7Cnm0n1
YB+SPbXGD6NGR8qDeRnyK79FvldbX5HLKhb3b2knYMdnuWxp0RZsPGtkGxVBewMY
ii0o/2RKx/GnavK6iSirM/qTQf7vNH3sO4j3GcKPskhvIACBakkFaE81g22YFjEL
ZekvFhlCeXHWSbG/nTXJQejgmMAvfXXiqAtqNUPlWPcXgK9wBVKdOBAvwk0FMadR
b8OBGQCRA9sjbCz3oybcZExawLEz1AyWfgELTDnrgh/+ub748wQZdFREEHZpPY6g
Mai2/2yuIMYO5AdSV8X1jAQ+pka96B+ij0nHyQZQanmx+ak38B5dTP9EyqKiRqup
IkKH1Fb740VbFaheW9LP7PR0p+Sd8vk9tltGY8TB6hbMnRm954nlV14ohoPvsiEQ
WO6R4ztKpZwmiIoxjF9D+7NCmrjYPfeGwOgIHYXD5BhrK+i8dTFWyQHB2eLiUzAS
Z+XZilmjKEmqQ2hSLngcailprzpM6qIgjq6tf8AECNa0V2cTG6zBz60LLQornEvj
N5/+uxgLrGmUQtz5Rp+cXB7g3bnN61WjKiNTHZuhwvRp4IhwVA0QFfUNdigboIod
jMvnJzq+e1n/q4SXxbUgfqNSjpCI8N4lmIV4RKa295W3qBkYwf1Ra//PlbAkuvZJ
qbuOun/0pSpzNxUFic2p62zbR2l9Yoq6VDF24dusUPwHMPkGmlkizVP4i6ZoCcc5
NGQoj6zDNUq5FEv6LUqoULnu/34tOo0EqzUxacgO9hMR6+a4TH0E3aGJRAO3CG2S
1AUMQ2EJwEPyfzfuLCx/+bbnY2s3G3mNMtzNUdVDVk/2zA6ZuQsLGwtKEz+XqDZV
L+/Bu6EpGFk8/tPfxkEl5LuUIj/mPh+vvqOdsqQo2J/qDWa9HLCgwA8DOvQczpW4
gvXvo6MjDTkBzCx2Zq0VQ7RWUDJYr973b2crvP92ulZiCor1mq3xhMumnWGmdblx
6qDd2eLEm/+TYckWId8QrMJCebk6nC8yVN36A6cYhlnoO64d365LOzVwHmoiB2xm
7Edx1HLla2iN3b1CJUYOVijzmiButD7LRnqNdQlxjlCykWReCq78+hDphAav4hmK
rTqGR6EOa1B6c8AtWWz5h/lghsSZIeMXERzRPAwZVYUKdBc/2nOmLBBbzrEP8r60
ClFYnFxn5PAsh2yJOjf/FBJFn/395ZXzou+NQhFCruTN3QY8TdS5KqdK98plyom1
2DbxWXTeuhnsEOa0Xghm8AiIMafvtBVbXJEM5AzMT2ToLtl9AijkkH6uUeJRrDfc
EKTUrvaczDV5Yi7KnVrvyeyEKgLk7Jx+gOe4agb2B61Gt4xMLLKp8RX6dOJ4G/Mb
7uJa9dKF13iHHQjEPSC+epAj561JNigOb3bm5dWX7HT/d4UP4arfepKSD02e6/Ds
Gm3S67Y1D9V7cFwfTxHgF3VRTSTV4jUKyB4mcjhjDzI/P68rZTjB6ltkv0hQDqbS
+gEr4iBlts4/MCs6Mpr0sRi7PQolauuB3rcnaqu4Pgg0LcZDPeh70Cnt/8+Uf1BJ
U50/CXGequx72gBilbFmY2m0zbF2NgZc9XwgduNOjm7rW6mRnfLJrpx0o84IplLD
YMlQiFgcJb6fYUsAL1F8Qyu3V8q5tsThgnZjaNbMDvwJbx7ofgNSoJc1m6s0V3DE
cje7tH1YHvO/BgTHNupGM62qdHJ1k5lyZrZjb+UohfvCEca8BxHV0CzAgLmzenb3
UmIbQsgLH0U56kGATgSDt//d0NZG8+2EaLcO7PMhcGB/17pLo+uAehSc+Ch2HDum
9ZyIEh3nI7Xfyu985XfbPNPqzAdmbTwWgM2izNcSV4eyMptL8Hps2ESq1qUz5vt+
qVQYWUxMHK3hd5M2j7aHT8BtdRKP4bQheQ2cDTlm/NRb9INl8F6FOrtd+XX2k0EK
Xep5tC6UuSvme33k14G2gbs89ejYgIAk3KtQJqha1izVXUXeacuSps20uQpz8b1q
MThW003eapPfvsDx+6/mtxZab3TMalUDLL8EZuArmdAnDlPuH8bTcP36Bbxp0M83
u8AFE1W44ku6BjJ8o/Gn9At8FxAj8YY7fNg48r5VqzS8erdOswjscfycJJeRC+5k
nalzYx/AQ1xVfkAqpEfIAFbdiWi6jX4FwPSOI7H/LwRMv+wqAgpOCRP1M9wdtHxg
mt4BIQ9D/6yIL7Kx/mLg3YAPy/HucXD1I3yJUENO5WqX1SWZd1tJq+UPSeQcQrmB
0lb0yLz1HBoTBQkdk7A6hdcC8KkIYfiebbyHzRLTQskUUDwm81OKyEJyjsGWopho
Nlmt1/phJc2+zmOoJfuqq7CHj31nKkvHzNGRAnl8ploOpwc4OagETqpPLUpsqgSt
884+E6d6dzk5S3rKptZT0+JdMmxuujBIglBs3fmI628J4oLRaKLInb2kK9bNLNq4
Q4hepdQu1RrvqBupjWSnUFhTBdOQMW12Mg+18loePdfxFemqkiY25N2zRzPdFiyx
td3lRSplIkXc8ENPuCCOtmcNJ1Z/8T6JQQgUmOjlhMbT0b+6H/eR01XEkGKxxTv7
xm/Gk9RH8mWduqsvhRfjKoxeNfzGY4ZQqVDu4IjzvBGAadH8Pho4S482Gzl6+Ouc
zMVWUkUPXZgygO+NKK8eBujS96V8zxlKDixtbn5k+FCYkR2F4c/CBAu0ZjAd6oqU
cPSAGSM+tC7G9wTaXEVbE4mxh6yaeVGbe4cfjwdCAUuDp2KnyDut++k8fifgGg74
/tCkRPE2InysecKv/Vqng+L7VqYAbw7gOnVd84cV9bX0mNNZ+OgaCgbm+aoOyir8
0qiSeWEsSgKhRmRwncN0iGXSfwaFqr7nLuRQxJX8GQLIhOtUZZcHHncYX2qMTMxb
zqAwFNpy6Q9Nc2Yz0lQFcRrW/lTxRjhta9YZxyWPcrpBJYGtV2NiKVUtbybbkTmO
p4kHjUcxUBB5HRxhclLkiBlHdafgTCo3YDVk2uHJwXc4tJhKLvpgMdEXRXleFyea
PwcJ2SKR4kRThoDgCfhUV6sCVKc+XhQOmi/DHDpaJtikLkA7HBFY9VQLw5dl7KnP
YMbxkpnq7+ah1K/J2HZeGEJn8O82fxgvWqG5SZN/QDlU0OS5dJZzHo6GqEMafQi9
tn4CeJ3Xb3R2oJupSLUusElFpqdtVYQM/2sCg8NbhW3PSMbZOLW31lNiAT218Dgm
j5sV5FfTyCohFGEvqe/5jb53FTgXirhJmJnIR3JpKOJi4y2Zq0j0N2WD+hyvu9EG
t+fPDZw4fWmJOSbTq/Ninb1dmu0+o9hz6xbz41S94NQSIbqJJdwQ72IEbWax1YMQ
kUYFrDF7Aa0VCLLP26pDdHlABtFXce9qFMPkisamhHfI/pqHPer1p+J6CfOFCnX2
Nqffr8fZXK14uuCwn73y09rLLti9yHecGEnXwyBKFIBBEZCamUw/rsPys8mJIdFr
fYrjgzKGY6N7dogPDlyJuFZY8mAFCCJQw4lKsVMU6d4CX3+ajB59nyo4QEnUgdf7
MD0fqZzO2blPXv1kuNV2OXf+bBw6+Fum3w1LWRNC8m2Ff+8LsYw5KvpUPK8oupNX
2Fs4H1GuXfTBIFAR298r/pIxvWd+edc7CKOwMtIr1yWLFl2sYOqBqfQn5BeFB0DL
AQWjx70cJYUpV86ErWvIX9qmAKn50Oe/7VFyhWTYnfYAlJQ93MRhtMfB88nIeovP
Uz1VePl6/+cjjOSmRNkJn/SbFw9wgCSOyho6UAQvEJV/iZGsvXwWkd7/Ot4kg3wz
CtXjZpr16saJxdVPdlmCcnQZvtIkjsBv2Rslwy94ge9JBHJrd7QlCtEG6+AK4wPV
zzkObPHgJku6SjENBbhPVMRcdzYw755EjtePj5Fh3N1MGj+QexQweTWL/jVvzhK6
vL2oh9u4nKkZzZgCqzdP/YC9tB1SCekBBAULaott6OTr0t1RoKIg5NmIqoPYEGe0
DqSkK5JRvaQ9Q4piR1PbHACXu6AEozCryH4ZsmdlN7Yti0eGkBBiq0a72G83D7ur
u5VSPk/wAdttD3XmqiXei7zsDZQGopkoseU0/Dk2QKtuhtNe/BrIX8izMHq4Q05e
Bnyzc65CjQ/Fh/3OnQcNEWBQFvWgSy7t5iBAve+mDt+yRatxdak2QcYfsZ0LvgdW
+E56FI+ibyXgxb2G6YiUSsuPbplLUfDeSauJMEueCycHZtvHnhrb6wCioct9/UDE
gSzLJHVOeChG1WbjGlEx9aw8HGBtl1/dfsH5h/JBdgxKCZqhsdMjBAzv2/DrShSm
jtjxINAde4gP8nDbLRsbLjVCWTqZ7Pyhj2IkYtgqwlzquERXVhdHCmWxSryrEIMK
o33CXYQ6UTw19HfJTc59BI8HuGFuPS5jkJMIVBebPz58OpYU9mJVFgTZPswsNx7Q
A83DYa4QyChHDME9j7ZOwQdybrvU/tvhbRRlFY95BHirA5dkk3RQxbL0P7h5Iwe7
wj2aoDpfyak7r1dVXTE+ssDMvVc84DxnPOVZ38mTMjwXGwCqbf8VYcvt1Y56SPxV
Gozj1O1m9aZ4WcRZCIXO+MGNLK3weN18pFuqhwTs9DDBRyreKCSiol+lGWmmP3sq
TtCz9LbkbD9og5e+rFHpXddlPjAJjYW1IcEfIRlaVxGI5XQt5wI/SPC1E6nVLO07
xlEXhQdJM4ioD6rCaupXIh3dPOjvWMes5KF2wHOsGtnwWXB7mKoECO20Qfu7BnPp
4BjdppcrKgIGBLZct7Vss3pLBBDPNnYCS2DIdWNv5y95u6P/ipEOerklTPES7/xH
nxwf5syAyhpMk+fjyy7P9rC2A0Gwudy45xMuTupVAiePCgp2L6np42lrNqbwz40w
rw9JlfeXolq+Sv7qOP/3GcMKBt0mk88AqA0LeMckr4pR9VRTkL5awlD5TqkvE262
+SHe+hthoNY/j47KjWiU5sJkac9i8RsoX8OTkhjCRZG5nKoApskz5s2oXhYEroKh
DzqZo370RDDMZE5CmiT/dIq7j5sGYv5ph/8n/i09a0JhlAUC/mMXNjZuQLhNg9vM
dqMqdGWzcuYM5hnfEL8vpQFi0ANDTxcfRlNzvGRoxtGl/hFS139NNHeCt/7N9VDW
KUVRFlrXP9FQ7Ti+FBmegHN7hMhEPfV7dA7aeIerJjHSI8dASfOHes2Pg630ONkU
KihfQ39mBwYGw5ccpce5xqza3+qsN38UJvV7uzrPsuOqZf6XNMJlGM5posOjCwG/
LdjAtYIedj6MYySdwY8MkHZ03+XVamkPFfTb5jHQvIHYRrGnvi5iLJYowuMvTCy4
bbnCpH8f65Jufi7r9bm5+EPpnRQ3JTvUhPb0SsgRHmn4VnUXNnX3mdTeb19J0gNu
M4BWMYH9j/XmXDvXqEvlgHrUs1VoNxwTRmcbRxvR3gPELIegV4Z+YIxN0uJExnYX
C2lMBzkwjZ/DtRAlEGSEVMJJzKqn/Vx6HgV5y7wbheMGH5WfAMkPUCUmfXOxofUg
WOJ3quARqcfwTiMhFxPCtSAOBZ5yF4hqB88CrfnAmmrBzR59P2wohK4DGhdb8WYD
sKqjkv6tR6oYTLySthRIr+A408OR0RFnXZcaJEHlygwo9J0Rq93aPDByk1U5R6zY
CC06t9G4CfAZAodFtUMh3ntd++bYeMwW5Z0Yp0D+mlVzn1L7mXJ+m5VleFjpHXza
+dDo1XjRK/4mVtr1vHjz59L/9ArlUAo3MzCmyEnGL+H6i0RBqQh6Plaz2VuDOWIK
siXWX2PW4VZpgugyEtnvcayFlZHWUsC5857vREKsPGwxjmGdigcufbtKlxc5Zd5v
SXmJinW660xd7X73CscRtpgHeWPoroco3aHOU7DMsHvsSElw2h/Ll00UdacHoqct
Syyw470shlGCnzdfqGtIW6LQgJ55Ty4NGqHO43DYt+r/RXCL0shfho6hvQL9H1cC
vJYjQklmqRw+e+NxJCKOZdHu6Uw5W9VafaVSL6ffFCgie5VE9ZrO0Wqz073506H+
16auvJVTr03/EWgyg3upF8aOpUpZjUHb2oZmYJKVIOqSHZ14UYXfdaYF4S6LKcdp
P6EP8vzm9JeKYl9LJOi74RKgUU2+mpfrG0MKTN4s2J8ipe2pDsLRXNm4aVMmplwV
YQKv2/bm584lAZ4JJnASCzKnKU2F8x8s7UrcqtDWxbry6MGGN2p1Kj+PJGoVkZfz
ZTPZOFeRT5HJvzv73q/Kyzv0hwYN1IDNxsYHVYvc1Y6gLx79GUSNCq+mNfKhAUff
39aLYjH+LQlutSRVJXxnPVUZKwcy4OSAvDF1Wh7j6/AyClrAYjqxuu96oLOwDB2a
cM18ImM9F6w1XZly1f2xOasykLXxajG2VKOPH1JF7rpZp+jkgIuZZ8/kJQrrkMkI
6LukyW73FnJ/VPNWdJ244gDJenNsxNlwYV5QFvKc1ablTXcEfOsHKyajyBhWVNrb
lNkju3ei2UoKaYXEW9urTQGjXkS1LxLkXnTOwEHVqXcHW/+Hi2p3hUyFjZTAShUR
ISbcm+7oPLPZIjkDAzW2jxXNX3HMB9yxc8u3S1vZzytCDaya/IlDg5Fsj53CWPhR
itEp+H5GqUazoGOpAz5hRcd/mS9gVcRHhb30I2L7QwkDy/nwTE1kZzlW9QjnDr0G
+f8o3YKbXDt0phMHm38ujOUJHbZQVISgLwEZuXjuPeYoHUHuSAY6WO7uHntg36FJ
zbKfRygBSKuRqoFv+atRcu1Tc/beLMBg52Zcrh5pZ36E50VZ5WYMwEnlPd51MIis
giXn+E3JdvNi4sibGpffW6/kKUr+tBEHFfFt2rhSnEflUA+rjItgjlGONF1Gi+gx
qvrtpKWko/tq/Fs0SH7sCpPs0YzYhzxFTDXppIuw1wAuIcxoFZHzfjMvg5ALJ2qg
00T/diqSPVjOrmapARJczx+gxS480bf9BWkX7t/QW0lmXtzyLZ+8SndrJeLkzuOD
OcnMiG5dUDH922ytle9nnYQeFHK7UO5W9l5GsGVJr1Be6QV3oUIt2Mamedur7WWi
spvTHNV+dwnCEHS7qVrXJktrTqMmtzCGN+C00LKPTwEjVQdw16+Ejz/tWx0hsFpS
DXAgS/KoHUy+Fru1gEfQlnR4Iw1BKoV4IlTU9JU0ScIZpI3wrjkpXvmIgovIu4dt
PgghXJ6qX4JE0CWNw0kKw2dVfWG8TLRbi+wp78ySBIhSJO7yEmYc2Q9ALrM/zA64
rmFWkxbaGd7SLFSkV09evA028Sr16NjqA27GVVa92k0g9xjFA2y3nbkCTXPlVGs+
8LsXUYplXKKb6KmRCiMKjWOH31/gXyEHSjR6Nmt9FTid4dmKaahgNHObWAH92NUF
DVJ/ueAG3zlBkOnD4+KC5oAA+1PVoK1gyTK9E7NY67AsJgsniaAe3QTg88h8GkBY
0mioPw6mPVwpCFTsK7kLt9arYXVN21h+kK42o77qYPuP8r68LBnkoju74zzjLGTC
uk9z2egizA72UkDe6T+CHRdHTC8DMsqRIYr2HD05Gma6x872lfYqEdR6E1ZOtDXn
4fsAi1xYqzQZ4LTIdBdYSzuI/Wr1yoq3kPgD1WYkW/UMFU6tSPVq3voBGt6crcn1
uuINvsGaVUIDbmm+XAweoXMI295D0q+cDw8oHa/3I5Wz9ZSHkFCYTnYHwjh+xb+r
mm7unyj2EiL1i6cIb/GKvHacAH+ve53SvVzGU+/iQW0gC0/sam/3eKEoKnVOTJKh
jh+gY3dMOwIaEjipwud5SXwxnfuXhBM4ck+Pl0gM/nyp7OjK4N3kOCTgMMnD3gHv
XlRtsupDjlqAM89BE0D19X9+6ztNS7pFC8QiGYCiubQ=
`protect END_PROTECTED
