`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYSV2uq8R1XxWCLpJlCD+eDegQjBjRrnXW3X4Ol+BLn70FYfZm0blWOBHw0UWPau
By6TKrFqeMkigEY9+QZXfiGIFwd3rjpFR0nVZPHhyPIP8Rh1yhSTuvWqRq3N8sKd
ijduyzMeVrjKx1/Nh5Nj8ZoSIq8BgXMj44ape5//97IEtAMk0If15uNV4WhYsuCg
50u3xOR++dYszqEGIkj1l8GAJDYmh+nB//YMJyaJ/TMUrz4l8Kss4g7xy25uh+hi
xeb0zJYBRNOTnDmJulOVHKGXwUR4e5M2vVYqXueAVW8XfeXOoYSMBXMIgwREIUhG
psaA99ZxWbD9gV35bEMPGvKeYPlq5/DdyrXCZ4Cb6HW+RG0DWq5n77i2Wq9QB8hJ
gWro5D9O7qEQPBRR1zx20ZUXAC7lSr/+XTyhsz3MkoXswpiF9u51Kq1xRAkew4/Q
eTPOVihN3DaruMEXhxiaxpvCNppqdd+jUuSrlEqQ7a2aYn1J8QYOdNvePpKyhw1x
gUPFxAR9demOgFHAaTTXjv6toDhhODZWXt3HexEOcn4BJBcUW0xVCD6JfPtsml+J
ov20G3imbc5LaCCH6TYasVEtApMMwlQe/zfgWKReO7KIlY2zUYO2CYrky6qdKhHS
E0EcHCBVwG/Ulf4XeqgNfaZQa2ae1QGP80cDtZeWlp7N4WfBWWetHzfEuKbCsSK2
XptMG4Q0Tk0n/SXSuCxa/ECJedOSKqblrpNk5Xi6GQpQDvl0ijSVMcUOyDYqod5w
5XqAMGgOiVaNLcYGKRdFzHcG9yGzs2jEz5KNmY/kFvhRuF9tHa0SvlufgcitUpHf
vKE+tve7qD3uin+7bkugyCqA7icmVUqbLW+LMHeHwYwdWgVqMGboLYYVXFzUANgw
oSCS39lB9/6J1uRaVRFzYvU/6Sw5u64vIgeStF6vUqD21XwlZZh7feZsNTMQcNI/
xFJJ1PWlRaRbNcQvDk6sBvgcr8bO3eo8i4FBxENJQqLEXYeAgZOjtZyed+LdKCUn
7rZlT1/NasmlBSPpoX+UWKN2RQGYyJOrpj7JXTEWWLA+xw5hv9q1sS2W/d6AEQwO
rkSc0NiWq9IgdbDvsfIrUdX8dCfI9fU4nqIjF0w+d+TvDwlW5cVFroJiYScNZOVq
+bNB4U6D4CQQmXbBzcVFoPmIrnxN+F4m1ueQYkX0sgRk3p5nGP7dTNcY3qj2q3+e
iM67xyfNBErTPm+z4kr4A7O4JyLD+C9u5B2LlMBbqzkx/ABCmJQ3PaVSHKJYLD6a
IT18iGkL5om5jm5UUZCLPl9gt1vjKh2mhoRwRMs9TMc+JUwNhpiPvflKn2HVbg36
AuvqJqdDuLLOaxbay328I4/BHBEixPtGPvtPxFJUjrVfSZbrp7GZVbe4hzlKrTbM
9VsKcHzvxid/XRKi0nr7/AEOAZwmznk9+DvNCfelw2oN9DORKR7fcK+Z+XAoGQbY
5mg4JBx+VkxKRNgyBonibFBu6AGl5XCHhftOffnBCtJKvpSb4giL7YgoOtwkQZCX
PlRdcCXHpBqdRDvYOPTLLjP5fhU9QvVfp504LoeZdxdj2pC4S49hcRJLsvfoM1aU
HMlYhLHLiUwhDrgi3J0Ij90SIqWpFLXAWKrDk1G1XAbpzLWFbxxtO1xLY3T7r5Kr
8FZzhk01lFvPUNDoUpdOI30wqY6kT/WZszYqs0Ran3P/eR32mAB2tu1WuN5NngKJ
quPQU5ssW6lrmZ3C+lz/0XywN/C52bJMo4qO+Ef+rWdo5qi+k0jI435B5jW+ph/P
L1XT5rYO5uwiwoyGLFXNHeU10ITDTA52ExZrZGXXuI9SkMrrudyE5bhfJMlflAdi
khwcWGFpHkk8jlnOcGWM4B0EkbbKAyPLIFFYXf64JanHUzPMbDNuCw6akeqbWsvV
1RAFk+40u5W/VV2vzb48oxWptHupjIFqWLnFq7qB6qoRYdHeqUk1q1XhN2srb0bh
Xo9lHt5Y+SihmWJ/7FcmAodKP8RJ3KJlHaoLoyapW7p7tb8Oh/lTGqgchSoISNHS
PJbXtIYLYLFK4NNsqbM3NQBP2zP9FHf8PRh8jeqD8XjPqLvyM+KcvB1GLjmcUKxo
nlje46t3+YdSyKuXhTCO5UuCo5EsVmhfxohMOFio4Nu7Zsr0/qHsDWzWTWHroI1e
QiLXmCrbJ3PoW3VR2GQNlBoD+zmi+fXyC24k89MLohU2k1eHBD7FQyvoc6c99Tal
M/hg0xBBW9koWq6IbJEDv0bIfoRS5uC0cqaSSiUQeAatyC+i65pePdPKuZ5kY0/q
hkL95EE0S5sU4bWBCHP/IK8lB7fopBIzqfnT/v8G6vIiurkqR6pw9ML7uM2HyRqC
Q1SnQY6eeOh1U2uki16fZyJytZMYzXJ+7w/ksrubgV5uOFwnxQ9HRtJoG2PwL2XO
nTVDKWWzQB7GopsPH1kAvw0T3xhfmV+6rDBaIR0hkt7NZ3AeMaprPb5vTnqyIlBD
MRYL90Q7OOTND48UZCj1gaV5ekWVx/LP2hqCxBMIFpDyH0KCgCx8QnaD+FH954uI
/5Zs7uCErHsexXrxZK/qzi7qGqzYN5Hu50uxts1ErtuqbDBzBccofD+0ng2F6CDo
Xs6SQ//X5CBStSYWMVeUuW7wJNzAuyc9KZie89n+7mMctXVrFRYgYEH0+neTYJ4W
cGcgZXYhetE1inO7NeKFJ34eAwxRtVnzQE+HuTJGKPMVyRDXSMGHN+RYLfQRpmyG
QiX1QDvfyph3qxCvjKxRpFhlDp08/DtEL+w9CJUM3Cc47/hle1o5m4CZq1w5/CSy
QkNr0HFxxzcaIrF0HHnKXVIIqTIQQ2T0Vd/s7JPkVNe2bxpeLesNDgJm3WDb2Xfi
UY/BLCM5g8HXZ3Ying8DP3UE1G6+a36WngOovhIqR7ESh3odBxFZOiEm1CqKmgYE
/BFyfckkLTQyCKk3l+fhGqIBVjSCtCkcWQjdLHaL+JWbrtxusbmWxEOAm0ACubiy
Z3pN/OH0MLTfPYAnXQsRs9+2xZrF+EWC0BSxFDGgB964XBCObPpwNfJaBhECbTGV
Lzp16YBb3kglEfN3K860J2+B1tAaWMSRRq9Txc75PWeFQq/p1cVyUk4HD6UNcMzb
iF6mWYtqN/Se+5v9kxis9MCO8ke3t+a/F1TdhG2P2Cu4qCscLkjIRHvU1m3gk4gV
+vAga3PV3nUqZlLSCokFPdXwHbvWR4qd9iIu7fiv0ujroL279MhF+EjEymajcNFe
VvsZsk/jWMqa5H86dtaIsRvLobCpntPGN7XjLOAeYMhnwjnwIARIL6st0lNBL9nz
9BZKhAAoMZYOxd5SuosTs0kpSIrGfUomXUnkm4/GkKchPTotk1BAyzpI2iUd/wPz
DE4QWfA7TwMGgJg11GpFkOmbP8nNRR5IJN3ii+waOBSGy4vezRa6abZ71eTsTi6K
Tld7PU6X9HtBDr1MAVimsJyt1X6EDwPxpYBuDYOXe3cVjrhdXtivph00TYVh4BJz
92TrKcUyHWvbCKTgOtoq8ShYo04Qcf4nsEYjbDUBJgeEDn72jbUzSeIqvwnQad4r
b4bFI4axXNNeyBAqa2MhttuKqQCUcp7zRCDYp6EA/NxpwZilpDunu/v5xrFKDEb7
uyu3ORChqDKnYqt589VwhWXUczZd8VMEcyDqEvmSHr0kLE+GhwfczBUjMKnnqD00
3dZ/QBBYT8BqelKT9vYCntOCbcpVLgLkrMFUhztavULzEXpnKh8hQXP0t4kW6xlk
+6yaoxATEE30KXa3FkABRZS02afpUHf2SUlPNQERJUf+4Ukc/QhxDDJNEpka5E8S
SksNNQVXfErqN9FHu/YCNPuU6G88ny2N6fa+LN3LRjtixRFk5f423jAdOwg+gZ51
PdEkQMU6fsd42tmmC5LeJwat1bigcu3hQ+VkteeSTqPwlFz0VIevl6+3N3LxiyfZ
GRdZS7eMHcxQgsPwwnY5jkPcfXlsB+t4Uc7z+cmkFVJG/vQy8uyYPtGnrdGWj/7o
d8EQfvOo3lWUDURMHk/k0Vq3UFa/ibbN2t023vqJkKTBbi+jni1OKvYYT5hAU060
3h5ba6fKWo1H+XsqO848Hybmx+UpLLKQXXnjTjl5BBOFxfJEBuR+78N9sneG/CUc
0P3CBqMNJOxYrqhborxW7u3kF/LLq8StE6DF9p0oAcLtHHG6nO7Zd7xnpqEARaxE
rikY0+uxhVE2UuaDqWVqUFfwpQJcRTmeEm0exjamCr3FIeZvvk5F2J/W1fRycWd5
gJF5XQeOMASuhgrOPdX1XR/F7+SFE9BVtJMyBgQZtDsoemIldKKJ5gXsG2s9EbLN
b3iOwt6pFX6FC7fpX6OetBlb1UnvsVgHEELBRVdLKV2roEpSMMJ95Jg+YPAp4glb
3CcKL8uO6HcVxhLnWA1cB8+1N12lIZiD/sDGiSPdgX8v6/hsIdgVBq/OvciWrjNF
10AUCnKl+dRG0bAawJYTar9R0s99tvBbuYi2F06xAhesxZ0DnhIRTONpVyBiT3Km
+TfEEjfXQ8YzGUckDkDQRiBLg7Nnash1CG227nhw1ypPhwBU8iA5ehxDySn9ORMJ
K0Aynugg9q9iZQQgvE20jAHpBOtS+s6NWm2Fw8oyZF9v8chK5JLHITQmwujEmUuB
L2XJHXxc1ZUVLg5mSHgAidGFEwQ14BxGJQQ2ldTCZAvx77fbYnIhkxAUUqElDb4i
ZWyqFzP/RcSSrW0ufccglnvu8f/ID1v5VPFldNUkm+K2jBJsaSu5rNx5+/6BXE3H
5NoCURxC86Ad2gjcbnW1Ntrz2MGl+RsDiygZv4PImfBvIwFId6s3H+u1gGkzUMqr
fLO88fMhDQ+RwVHt/wICYqDPGCDDw3SjCb7aw/EyiLBi00l5UGjohXTpcdjUlwNC
BFw3B3ZMocFoY2H8/F92IUWIAUC1DZKaJOnkohfxApvIKfFrFHXxbiILnrpKUtOh
CsPHORfHq+3L1gZI9ttZLgzOm5mroUolDfxSNBF9JPQAUoCO5jFYNTE/wx49iEvM
NJHu65eJbdvcft85a7w3PDFjaHoMNtlAcWpTAEGJ94hFD3j7FgLB1ifz/AT8odC/
2Caz7EASFomFoB/Ct4KVP6XVaIJ5iW79VrpKEJZFbxpWyLkWPy7ugFFjnpQEhxw/
nNZDSxwu/d0dcnrtlh1WDU4IfXonfADtgFB+ObkW+hrw12ZPnqq3pmfZOIgoIoqe
+FHwt2MK9VWJdqzEFIpTLPu8gou6kxDVNsIRXq1M6gYdPqU+SYJTtcbUN4DB1aoi
MI17iJEeVU6YWYHjH8Jan3fRyrXq1S/dYsExiYoNv7GcR6zTieg9KPIJwsEMIA0M
3QkqV4n/uHBpCq/vqaGQEIcT5FQ/0+5Uuu5gIS5YP5w9p933VegXR6/5FX+69lwp
JBDIzPTKt3uB8ir2gzsvnOZ21llYk/vPRnhhAJaDkqlQhFWUNvxPjPmFM3qZsEhh
/ogmLTqEFXPSX4effcH2cVQEJRqzpaA+nYlHSgMLJRLPBIYdwqdwLUs10sgSFAK1
r1G6drwvTju2g5e3v4CODEdp0ZBoHkXI6XjzFUVsR8m5lQ0kyw8MxoUJ3eiX5FDe
rQ/OK47M2/9yF+v8a/ypPKuw5+n7fvmTlfT4csdo+oaauMEHifkjhTK9yvyQvZyY
UECsD316xkGSq0E7wvJkQ0PE7HBQPN4KNAGu+Iuk9PnPyo5n6ua9PvbLocTdu4qP
Y57NSUpCoZOhGMdElkLhK83Hyn2GVeQrT/x0EzHqV9Nmz20oGLneKEqn5Ad9h9qi
nqPjpx6ZluoVmhXF6jNlAMp9f90smaNw6pZ1H0p/91bQzUKGExJNDcRW2uKwRO9G
qMDJ9i62DpQ2BtkE6nxAFuuv2CCf/Eq8B3Qfx8SMJUk65XHvd+fumlQaCZGWfFCY
tyqMTxPLLXyZnowoRgUA9udBaXxwzwaErEqEOlN1BxUDWfkwHxkyMR5riDPEl81t
mLVHkkmP4uSZa5m9HpTRaS9dLZWPq+AX44BqaQY9l0rn5bDYMATyBuiqHNve5sZr
K3s8VuHDWfR5jMq00xR1Ivx0TnKUy3zK6jayIlU1dENPhqJdFRqkwEQnh1cgjOhL
a+Q62X8EARS+Qn4c14idI26Gv0M8rXQ6hi9vvxoP++aAjN7lkyQKv2Slow2m0+Ql
/Y3Vd4wCbTeeeqcsXaEbexATXHkxRCi8pqRxLBVtF+/niQPkgRMPbg/6lawrJAt/
bIU0PPoZNoYoPpubAKohvEBkVPonBiOigOCWagf2j4lF7RxeU/eyT0SJ5ua1fSPH
VHvfZNbXhq1aTLy6IlIxpTyCqUiRg5k55qPF/TGXoMLD5NsReqGZxa/eemNDzTz5
lZoV6U1BjZXG7c4YJW4LZWMe3cGypci2YydbxTkWkMz6Jb1seHWi+6A9ST0xgVcE
8Jz0Quh7GhdJU2mEBeZxGt8zei7S1QObNa5CQT0usbdcqABp/fPTy5QSUiVJbf/T
rh7PXm6q1DDTKW46dLif1L6Mx3rkbyrYbwGRu4/LOy4gQkbcTN76Lpky0A1Lsld9
q8eDq0ViKlTC/AHp8gQ1Z4Lu3qBoj/qhakqRnXUK9eJ4Az1R2AQ7l9IbzNhcC+/4
yT5G7denqAr3dsgkoBBoGNzAc8tKs/gnta9TCqyYWgD2gQVrJnR1qtsVZm5xqaY2
TedHK7inya38Oe7hkgXCj8/cDOvmT1ROIXL76QdQKQcPRUw7UWMm3Xmh0Ajr1ewg
UEm7iH5Kwes7Iy175krur9YZHrs7tQjtOj3Q8C0lxq/KZ0PA8RVRWZdn2aibA1HA
VU6VW/7yhn+WRvrqI13uPTkOEY6YU5aMMvG2ySqHkwsumdNHaZd+mCJucguVuO2C
EXbvUMsstfTkyjrQ8B9MC/8pcH6mWxAn76os5JVXFq71f/lovJVFJXgu0+zPrTL0
s7z0ojCFKtD1pi7Ibqan0rIlovICHosx29NxVboj6fuu/SlgXq+O61ht4RtOq1v1
QHu0T6bTBuJ97Vj2RKS1IzaQVDijGIddxPKPYNjClyIfvvMPr37bxcY8KE9TBTlV
3Ymh2PsVbjsD5NHpgUuoiFXY1vlelxycwTfZFa4iZp8/6ooZvBX/kX2BkzHiYByJ
RIYUEfreQX2UJwHVoQM/1pEnXuSvlRsgZq7Bk3KAsSwZ9zNzC/0yRpxZ2TTAELJm
0aVoJfEvcLWxkDlkrarb5k4Lj6D+f8W659yrxmWV7vJdPP4YYbUSJQ9c0MYYEjLV
X8kmpwjl9ufRdUMbYHDPz8Kc8vbU+QrPw4Hi2zZoCwsRh4R5hi8JXzheD4wOdJpx
ubSk86E+sQUrJaoc7/NFsh4Xg76rd3uLXL73EKdXe/Hb/yMCCa/iqUaJVoft80AB
s6FRApRHWLnYufwwNg/vG3TQ9d1ZHjOlN7SuMqNAgVeDx4VTcFrWAZDRcHHBLQpk
Y9kXT5TyOXF5xi461+yLIKK9kSmuvNJArxy/cg/5nSO5jZJrhmMWB16+p5tu6kt0
6WdOrCnDJ6StMwaadPGNFZPondXFSrFxlAXqKL2QNJGYydYXuQeEeenGoGeA2xx2
RNtTcsySn+/RWIRWW4ieScYPrAnspkOPrv+CisDN8JqHcuBgJZMuuhcGvovCASfk
GzMGVrrRWbF4rSKC8LC3hYbel8cR/ZyiEI0horcNjW/ZFXp2bjgNko+E4PvTmf91
+PxFrpKwfKar6xPD0ROWZE/JJEYdkFZjBI//KGgdBbYNy9IBiYE1daMgcuxJPI1A
GtA/iGA4nCRNNZ/lZvOMmKaL4Qctl2aqJz/QvtGE5SOKQ4BQpPT++fuBOcbbqU6m
dZFISWBcJ65em88VPjhGeiuStCZtsW5KsaBzuzgzfS00MlL2orNVw480xD2a5qHD
8qgA7jv97Ei+skHV5WXaqLrOW+EntFSEDchwaGIJeN4f5J4PZacfeMhnlf8kE+ZB
mQbbPB2b/42BJuZ5jd94JO5is9WFc/4bVwlKgf74m5tiHJJwf5niDzEq3OYn1RT2
hwDJa4rp1A+BlCWsI6wZb6J8uJAz06/Es7K7ia5FiQ52g9s2fZB9xKv9usMoPTBI
/Z4uFooSLbkXm3JHiFb24UzJRjkPrS/XBPe0drZSk5rn2oJzPyk6EBZhyo7rHq7u
RReb20Az7hJ6E3U4L/hGwjdDL7rKK7ImXtXK01xEiyYkO1QkU18DK2JDmXcgl4rB
2jABK1b6qR1IIzVAeEl7dNUgQYT5yVpL/30JJuqaUWdS5U+YjTf+16sjP7Nuv+kR
quWeEEKnaWruUg1VNAHJGT7KNcImUbSA+uTVcDEP75eOGIygf73pjXjDD5uOpwxb
RLGT3ePEiG/XjxNifvnvjfXPQOHUn7G/dOL2Io4muAzEjzrxrbJeyl55Rwnv+z34
f19ZZEsar0Dt0dZTZxOHA8TEOpBPbihymCBMa4n+w9vZ5wHflIxwkbSJ4c6Y8Tkg
Xmujap068nbTNA/1BOBoXZ9/1oyc0j8qf+42/mcEa0drcX5IddrBGvc78ivK+QIW
ENQuvLD0QbJkrKAcgLt4na8wM4AkAwxg7r9hlg/9yAMkDSzWu/KE7et7elhg2m96
UKk/rM5EYei3amkXgHZRmks5X8bl/fbbpy5Bu2JQjA9M3Wbrx18d0ZDyQp8blqUy
OlSkNRE+422PYjd74mmH0TYp8ITkpQHdy8/hkptB2UyF52HV/2NCYyC3FYEK4WcJ
L6n3bD+W6NMozV5Fsgomfvbf+ZS/aRXjnP+dGm67tYPMyupkhLoMoYlzL7mDynic
/dJL6miAt/wBzhYzH/Xdnyv6tSnd4685qnU7mZmMoKmOL7FJvcURkN+u8GPTawBJ
0IwtiQCG2kLburSw4HugXQiv2nIy3Xa4he7ZOqnDwSE=
`protect END_PROTECTED
