`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IZtKmb+yddIwniNVB+ZRt/98n0L9mWdooVNrPkPvuri6CRl+zR+bJEnLnX5Tyni
MkzHH4jonR4h8EjRKAooYTcvOsc1LVWvZbPY1e9ha/mV0+LHsFq8Tv4KIi97+KC2
9oWFpjC7airoaNhf/RAit4r+JHn6ofFEdVJyUwAi1tiJBJuGv6Ng7BZ0BbtWzvwN
33zu+ZXhJUcMuqi8BTli5HsRCWtkWiDUWwIBt/A0sLihOpt/VZITPbgFS4E4Mmdn
ZgBHJmI8iOtrKz2yTUHs3t80cyYmJbb8PS/Xowi22A7C26y/kkZGajD14df67PXi
WSjfxZM9LR3dJczjebKWnSfhi2rnlV1TPveZcQpdO/qWT+OKhhTYGEHbVoO71bhZ
V0zR9wtMeMa/HjwtnX4WgYaPwBGObT+LwOmTEVx64SD0jdzzox5/BqQaXhAjaQeC
4Ch62ej74zg8GegNqtrb2W9LnQTvTvtjvrUJF9jNUbgehOYWLasZcWGqXw/cmuP1
Q/0EnVI/dmyVRCQGgXq0aGucLwVZXoJ5e+MqwxlFO9wIGGjJRMXPXmcb6ZvrmioN
hFhb6Z+9ybNEUTup/cnf4EaVTwnsXyUIyrXpOo4+LkyEzH5ajKKNvH4f9+HXSmpc
wC9ElTHHeELmWewQwY7hNYv2LUxGlCTa8UcXxftEleqBacxsMqnuqWNruKSja1yq
35LR6nbrIlSSTLGFjgU3ww77i58drxzwA/rpJ2ycPwjGfWz4RogvlTFYZo5JBx+s
5vbK4VndwHvsLj0Xp5FMl5BU3fgc9VCkkGR9WHPTuD0EJ+uC7CWu0ureHbnBrckN
OLI94HNIm3BSK4v/16n4FIsYiFocHvMgapskgGD11ABWyczvcak8gGlpJn1YFmLV
Bpn4ZV/I19T53W3l/ct8AREzybuzfKOVuXxW5YzqtJA4BQD1UsXOiNkc2qdGgHG9
NHm/uVg9LCqrtotuX3KgjZ28NvutdP/DyGnq8xk5MoNWlpHRpGlidDA7QptmGgSK
3VcSFL86vGBcJ7WYJ25YtH2K/LZ8pZ1nYuDVWxg6IGNSxRAhoPBVHX6OYwFgg056
4Jq61MAnxrwbj4pKxrmnFhINq/KEXiJ7ijSiQCHsYlD/c4q/2cJft4G6uTHncnh0
9EZYtAsT1Pcu51nVGgs+Hw27hWzCEQ/12tboa12Ps896jixLuGrNpawtjfgKuWR8
h1RdJFRdjfF70mMcPownIS5/1gI6yIDZ07fhCXBd2U8=
`protect END_PROTECTED
