library verilog;
use verilog.vl_types.all;
entity decod2_4_vlg_vec_tst is
end decod2_4_vlg_vec_tst;
