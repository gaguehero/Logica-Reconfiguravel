`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5eTrhQkxVhtqNgQZar2gjhlVv2nb5nbI4i0poytrutCkehs+sZfblg0KIwSd/dR
0V3Y0ftTr+deh65eX3r0xyi9VLVhZqKTlgNIm0c7Dfqedoh7BRLleS991khQIHI0
pcaEe5JL+f+TdxwRa/BRVL7u52lJVz04S3yd9F0fHX7IzRA2boj/AL9L9SVWTowh
u8rF/S7mfTNLbPtVZ3uF2p9kr5owOV5zFbz+hVHEtesYnFvL5Jlw+UAsEf5BK+Am
rn9sM93/3nSu29Ql4zNuw6EiJJJlcn7qus2BJrPRkLHAUDFerM8xpfgMJsHbyYv6
VtAhRO5+IcRUKLXPAQ2BYyIqgCglsDRl6IqvdcQNIE1j0LwILN4P2jDZ9uDHzXzj
xHHyzqQbZ1oOySreCbIHfvI9Zh0+k6YuFMtRkc5ru39Dtyatj1s3MJrJikg4T361
UkBgqvTz2p/ro1/WCiU2fsK5a/bSTltfGPakCw8U5+QT/qOj/kou0OhIcP8IpSw1
ojkZdB9snGD+7+cd0pPiEskaH9WEbGOANo+simVtexTVaPdGyyN/VJ4C35x2Tlnt
LyiMwhy3xk73tJLxzKaza2xowDuVUaSqQ4nBJ875KtIkQEEDyGRNcnUXJ3aHzCVp
2y+oJqiftdUEfy6KyWay0vWQAsgfyXSN3vJ2n3RdABtEWyXy9av91y8p8s31NDAx
k7nJgfaVep6NB1hG9xpjPFyp1dLbHle+L1KAipNQXKR39ORTh6ZSOMun3jQuRbmO
OFoaWeSSiHOGWgCF8VCYVQnmE+NbM0LoQXknohL5A2oYOvJU8Wq0Sh6/OFIhmfOF
EvssiQhUh0g1NsZPvWRiYOUbOjjRQ7azLo+gv3MtVMJWgkAJRVlebWVxcn7Vtf7u
JsDr8pLh/h3m4hN149HXX01m0ZzRuDksbjOrZskKNA7c1h/dp3fiNjLAzBoeuW1e
cFDkoBen7wGF0wfpXa4xK79Ojey2jQV9Gv0NSJcayyqx7HotJfuRtycJyLS+++fc
cci0+Ch2blxC1rYklleD6KTt0faG1Kmajl0j1stIwz4ZxtX7tW3eUfS3IxefSWyX
k918gBZ5Iqb7+iyOuesvf6+LhEVU/nz/xlmXOjlZCGjfkjOqzSGTxT8hZpcx0eNj
IkgS7XKAnl+xX8pQe8oANtESLbap+tFkloi77WsmrwzhF4JG7NacBn89GQAJl/XT
XMud4mo+jhA1Gbf6plIrcZEL7TtS5rV/oXI0XKpKwN0TmDlyKo6muvXHSmaF/J79
JwWhcRyCKzm26qqQkYrmUs45EQKya3PtUHG2pZfNLzuijJB69B9HnZSqOTsxbsP2
p/a/um+ElX80N1ZVIwJYW/ZIVsZEanvqbn6pnwcOetQF/z3jhL9Ux2KJrkole8yw
+3qQppOHMZQssBFPLn4W7zFO2WukJe0NYvHfTsRbBYjZZGJu2DIbafCoAI0doF7z
t9F3bk8ppe9bgGW3Y0T4BQavMzNB6cUna3V1wAe21MlB8QLc5GZLGyq0qOmiFI7a
gLbNGLedyh7SDOL1Jt5b8Hd68qbeO6Q2turxx4CmX2nSR2dC5jGLzA854HaR6ASS
OkJ30WV5K/uJ9CJ1ueQ7Y9plBf/qsIqVj7dMQBgUMInvJsWHrH84g2h9bb/7ArUd
eA+NoMxvO395xJgjZ05lWztP/LhdgRhy5rNw7OYk55hDnS7tmPWcv8FT5yc5ixLv
kTM8+WDkg4ErWYZyNOe2h6MzD0VIlhXMga8sIiRKCcrljVWLf0Mi8ALrHIJ+AUwi
zwEwcS3FESNJ0+O5wZlbSbvAOLEL32wkuPuTGPtbhjXogjVEF7Y52YSHdYJz5GET
GhxvOYxxrr1UYqrXeBc7FmnbFf/CHgFka1p+OJ1Md9DeJlXy4rDw2I44dxeYDzOw
MtjjgO5lEL/ZsQ2ntedFrRBFbTakliPD1sPDN7bfSOI0fxHjvKxXK7DIX4tNJfXw
aJ/OxNHFMKDpi3Lw7dziayJnAE4Ejj9k6nUTt/QyaFDsVK+QMOQEsz1Guc3k9JKh
`protect END_PROTECTED
