`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kMY8MEox3KkDicgUETghtEGef33ez1px7lY6WjuMu4PFdgOk9/Ss3ZPXte1r68rd
xFMOol4mSeT6THvQ7SEiOmhu2KRG6mdGqZT9UsPWPvHdt6seXDlxpmrGxDHkgxiT
kkmJdfOTckUOJyH9GKljgn+nG43Vm8PKPmfEd8t1xXk+AZwJTfZxkhAwGCsoJ0m9
gGgxodvZ3Mb6PoLtU9nvgzekZsID4NbbtGSrxut/bPPzNGB/ao+b4F/t0rwZDwrG
5RFwqfrpY+W22KVVKoQL1vNsJxEkvF7pzyPrDxSkF0pWJHhDex9qQKoinHdqvWwp
vrOZWto0FXsSenduDbfV+gSBJXeD3Fen0IpbBpvsmqst6tzwAn2X4qIdfKi3XS5f
6jwbhNC9lJJFf9GOJZydgqY+sIAupGFb7FZkcBMWYG8DWWaQrVFuvyiH29slgkxI
aUxJGsGC7VGXNJ2+id9B+ZmntHwfsKhVJC58DJ4O2JAE8c48RDnLMbvZRkawTYzS
jowlaMpq5Yy6OigGS2KZgp8qpO3yCZWOOiGJKO8WzaBjD8wSinoKx0gNAD6qEvq8
yea2uxYTExGSJVLFe9ENE7UsDyDzZGJAypdQWwAZI/bZnqoxzAp7msUtGffV/B+H
S6ccA6neY6HKGVyVOp6N3ggjjnB4tumRx8ZFA6ks0G0+XAYLdD2JmTOmGYjvpHr+
63vVCr8aaOEC+ONo6I3Y4YnTzAbNO5kw16QatmUj9xg+c8bjVn0rI1Yeg7kEF9es
MBSwvtmVgUgtRxdW+6mmhQdWNZviXWDIUr+J4vCMYdL4nJD+Z5xsePtapCma4R9X
wnAE+Wj+VCQZ/DR3j2J4tjxfGG0FLybuoMO3t1ZYS5zO1d2PMZbM8qLOxOLbue45
YjLyuEnBsNeIwaBCwWJv35mor+aWdbKa2zFS6QZHhaG3BV3hvCPVhi4bWE92rmGG
MevvtH9KHWA21OBYW14sK/DK/udBPZcG5EZq4MmYS2pGAtnnJhcUQzap93ffJfX/
7PDz7GbfZIrOpjIwrrEiMrzi9CwD1YEwfruFjKxLCni/6i5cSh33KwzSkyvDlh+g
nJS/5MyhmAP5UO/5Tz0yX4GyT8V881obc5ffZv7nL60haEGUZce58IOQicChFJOg
LGcedVMee6kC5ST9jTFJL1Fn4h/y0ZHFUoDEcSaKyFv2XEq4pqQ82Gqvj3cCuFiG
gcX2l6cnq5AdTnnSbAqTokSw4UY18zQnA0cFg5Ux689FeD52s17cw2bugz1K5EL7
yZbEd+LsD6CTvGz2vb+ydk7m4N20jt97IitFImiJhzVD5Zb0Mno26+Z9FXj8zf1/
KZuGRpC1x10J1Seu8ByVnVfVi+pqifmMmW1IE+inzLxJ2lSv1GpGb4OZpQKAdiNW
G9hrg77uwtd9Nr4CxCy1RIngyQ33CDALAG7v5fOLPEWGNa+zlIC18HYbj8LthoIN
BKP8n2yZsV8gKe9Y8tuACvD4qwDtabAb4UCPfSjWG2/dkUSeOgUZxuAKc5mtbfL7
6Y6CxD8WLccqJP7ZidzSXhpJeKjhYYptyS/9d1qBCvhPTrA+J5Jh5YswRAdTraXB
Ot+Cj6GIlotwu2R9X3KCESKtoefLaRZ0wXM5gF+ZxQACaBxvCJSwllUXEO7Rlabw
ul5LAFCwmp17FoyYGMTwEJAhn4jO3qkj5qXgsK1KFJcrIHiLymyo33buyIAGS7+p
Ii22jbKHxygBRA2sSGGvrWCO+uqZKaByuaNB2dGTJRvAvqBJAoKGhruGsGAA54dM
LE594SxRrhCS8LV8VFhRGjUtOpindOR6mXBJnQpRh9rSRe1RohAA8wRi0J4BFxw5
DmPeYa6OIqmvKpdlJl+IH5s35FzHz1dQtC07IxrplAAY5td4cXJ+c6y9GC/BrEAt
ZR5Zb72xVNA+sZo3jX1+sDlVzoaE/P9DHWQLnRDVs9UT8WPorWgYVFMQzYeXbd4d
gKBMBQ6yJyXAzUy3qS5fs+WXxm29UsZvAYL7ICS41MMv7Px2MGkqf0jwIYjIxaSk
VJlaMMkGsh/9yKyMAs0Vasyc6b0hn0QtGI9w5YQvnOz90EybPtjx5fEpRHF5V76d
+E9BmqKtWprCeBJSB3o0XYZCm0eZZKbpVC8rurOck7LYNihz+j4HoVx82GeyE/3v
udIUySKLh7RMqgEKeYdiRBWKiU7moJGsPBj6JpbSgAK+6bwMVKiBDEITZDaiiXvl
pIKHM7pUHGN9aUD9DscNQkM/iUgVeDjdW2DQ3jEQq46dwPh79CINs3XotfBl3ilP
GcUKdS5HUEGBOJLTpmyKvD5IKqzDxFao1Cn1haZkotMyhrv09xh10bZ7bgr8yL5Y
iRok2iJsqFUJpZYNQ9f+g4rqIhULORtCg3tul33m9XOAfyc6opPIheyBk7UtJwsH
xWPEiIAP6SMlyZJ0Z3vOYtq25MsHzsW2gu2qTCM1FKet74VLa8/WLtvClpuHTLwQ
KiwlqZhoOnB3tu/sXI0dwmzd1RrefgYqo+zKlnleQjj8CXOUF3B3X1pn3OBnduKD
N7xtkcpWRSPt14cwiXlcfLM5BybTHFNSLYmfJ52qbbFWttGv+ut5YTWJbenN/Zz1
766NUZXnuEM82955J8SWDCQ9NVtXGnMsWl4WXbWqsd/GSSW2vvIJOMQJVQnkQAgN
QBn+bv5wHGJ6V0ocYeLWlgvwdO5Wm3W6hPIG7XCifWi0H/8GciDROm8WVAAB3HRX
Ft4go3Sy8Zyf7MlfYJPEt/4a4xuuauVyiNHsUNoMjH5ImiXbJQ3XkTb3xqkXQdnb
CXtbSnIKPuuFk6QsumCBWWimrs82ZlL8u4+Gv2IJv4FYjLyhU089mtaX2EDweWSI
qd8j2T0+2LUTJHOxWHVLdsLHikWlm5bjtO8X0iaXu+oCvNjv0BPsgMDvd3HT9PZo
hCdK0JSbWI1bIZ7OxSSHC0aAksWcaQkOpT9Evbio+xKvgJQVYfm6uBDReEgZgeU0
U/kzOX/SZYr6aMX/b1qyeeA2LRPZWF8bonu/WhSGQSBiN4A5KL7PSGdiPhpfcRb7
lc2Qg1Lfp5+aPKB/oVME5fuHewBG+mOp87DJNz6uhBxBiI2lRHPQGndxygsSnW/9
lu8XBWoZ1NKELR/mJrbVvxRmLgik5HmBlYNI1aquJQmxSkg/mjYxvQ551F/qS3+8
8FCU5p+d7cy+rn/wiQu2wG9bXYWKr2rhbesUECrBnpoVbffTcVTPWlXsmj+rBSUC
bKv1azCgMA3X9isnwHXQDmUTf8hpL/QaYG0eCRu38QTlxWeH6NuZ/JscY6bvL5I8
g6egAj4aZSgnGOaB6++XR2tv5H0r5wpxWGKR0ar457VACsUNFWk92IYLBaXCRexr
jzBPy7EhPtJMOwAE/RZC19Sz4f6HyMd/B2iIgVQF/u7I9uE/q2JmkdQ6CUnk+uQQ
Ue2t2JEKDcP8dV3w+IFO1muuYlLsuRd070jQWtfMiPeTxLVBOHOdMKGw+0bkAjik
34GvYe+kF4M5qageWcDNXlWDpVHGii33clJDbO8deROW72QQ0b9/s9TKxD+P5AL6
YdhedLgfMVaVWLumaFFHFbe8uKBNlaWs61w8YyyPGXaatHtAEjOZRE5B83Cudelf
h5h+mr/JYf+3mId0rGXEYrg1Z73wD8RjQc1UpeEReJMttIQGhOR6Xg42NMlEuKji
kDECuURGfEcIVrkda1uW5LUXDfCEuXk+U/s3VrOon2X/OrmUS3Bx7gsoyS0cSzNO
HsA2NZUyMEpwUMG4K4LbiYvTgl2TF4PgJCysErubmjAg+vARrp19m9OYW1jocImL
FoYNc1VqsdOEtrrgDhgWTNxBfDZ+RowPaowF7UwFPPtIB8J0GNJ0sEtTen9U8C1D
peERkOxWZ0aUmXE+1hdMCu8rfVA0OwUPnWChMC5G4Fo+es/E38QyMe5fe2WJBbEb
bBHsc1jqwC49It4oxPY2oGtBQDymP8UXSXhgusjGXmNbVFcsgFc5cuiab/y1fAMA
rxsyfmgZo1VjdUnjFw1tPLUfxtnkJi5xTbvuSLTGIAbEM1c8EY5PZlPB1FicQPe1
IJWLwo9iGdkSMgRvfGIXefrQtmGh2Odtfga9ehugIa30ji9EUZcF+/Z67LCGcEpl
TnUTNFr6cMUUKFJAj+v9fuGZrW+vT17Dm6SxiI48Tn9YF8Hb2cJPhaRurT5JYh5B
savN4fPS+WoAHrVN7tLUrAgAOEfXLxBycstKltGUQESv/kd9CYHphUTw8n6ykH1F
xz9hN5pJO20iELZe56YzrCuosDOGS3F7KyotXbAtqvJnd0NyHd2IeMhQ2G+k+M3I
4LeJuDQaUoU0Uhst+6tVzITV7XzlNI5q9aMEUwZb+Oe13zUoiaN9b7Iswbr4c6Qk
d7v3kXpgenaVSbWdcGzbClM4ydZRWs9MuRxlAcqUubTkmiiFtbAe8XS0EeTkCom7
47vesV9Xj7WfILxh/UehRv8yjuTAKsHerkfxg/T3zGPkTsCQZkKhS29a/ihsHvJv
HPSuK+VfjNrSMEMpMiiT8dxO0Ag8ygFvid2AD82Nv3gwj/6E5rYXTKmDjzu2++6A
A2q5Vo29n9htBoeYjFy82MnugZ6NKQrBg5uFcGxx5QkIbPZVy2fN/ewmKYTWkPjS
9Bys4n411FOG+TeqAHEH+mTlTs7nGzyrKF50cvkRq3j4SXhsyRj0Yrbapp8yOkwj
gQ0Sb+4YNCZ5/JzBoV/dw+G+W0vBhdwTyDsZkUOiwW4r8/Ls2lG+UzAHfdJQIUDm
wPi8w7IR6dNsA8qMVMysmC+bZ/KDwHL2aDd6dshMRwCH6oxq3rU8K/ssx9+utSfe
V3SQNjPqNrsKueUMZhJnbebtNpHheCw9DWcJSJ6hJdUw74VhoySu85/cu8k3k0BW
pcZypZlH8tqsD2Np+fyhS2HMT6rfnXvBiQoJtYFA70J56m+mPKsupLCYsYtpwVLx
EeQXRXQmGDMLCpVh4oywuaGiAngfCkCitKo3HlkPN5HKV1QLedGzluAVW9AQp06x
H62DQOz1lFX+BGdPFqaMM4GjIiIAlPorsrgb1xfcuYOqJl0q78mxX3QoRVa5eVLU
K8MAg6Qm10OnJNRpdwH8lRNtyLymcTVdzD81VAYNfUumWP+CSkMA53kAa2F6UEd8
o74QMrTGdP8EYa2hB8s56/oTtWaMOIyw38ao7G1FrDbvdgzsUz0EGvmn9PSS4Gc0
25BCn/+9oy8ufo1M1+FqugiqtoOU2YGpBjKCE8NyVv3LuxCVJ/IcJQkL6uR6Ca2Y
lDq6NNa/ydgEmeZa8Ro4EvctuCMBD1ldWktt1EUqq9zHI7lXDpjmWp+qUzHo3ucm
9z/Ap7X7CbDXY2UcbSnaBF93TU9IMm0/5JyCpOPLWZcOOdGuukoEc42BzHxCXZLW
R8HxbkTzkXYfbWGBbU2ASj4ZIorxnynUZo3vlYzD2AgAf3YSGrBjP8+cUnIdJsOw
VXstCff5hMLBJT1HcKWLJ8LPiGGWo2GG8I4ptZuphexgCyJyFqeiI+P5IH/4vwAV
/ldbP2tAhtAYIuU5sES20nAOA/jOW4eaMA138id0LrfdeLVzuFh/81efd5AkG6uZ
c8o/YWTgs8+xHtYvgWBhLKzuUU2zhK0quiteYFvY6CXHNCRUYzza5Aw9A+uaTkmF
`protect END_PROTECTED
