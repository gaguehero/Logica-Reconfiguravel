`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7u0y1OPGzsJ0G9ncPkHChs475Q2E6mwtFYqmNiEBwaQwablCkBf+wvyJjW+bfim
ub0OJP55qvnnFs97obgYVnh9XQ9PPpA5UZjTyY60umDbw3TynqCSW1jfDbEVed5f
cu5WPdA3Dk/onWRP1jLRhtIVU2ldiIn2CQcEDVR+2O1Pt1ucQB1l5mUDjuYS3noJ
k07NAVPISuJ3Q5zKyu/r9NR5sp+muWhSSWwZpg3v5m3S+92sTNaWQmTcf9oPKNan
fyouVZ9nW67g1IA9Uhba7sOw4JXvkUJSXw7n72FKNtsgs7m/Zlf7jr1DJgdMNu/x
1y8LFZ7bppT8hylMRXjKq9AhrgpIWGNfAyR0vPA3rZqRyDBAGE+8hJJrnVtWOLIS
PPq3YGt75uv0dFJpCIOd/oFQ1lo2kW37An62ajG4TeG0ag5Ttr8TJF0Bad5J5H+C
tuUReev1zfLxFessvwu4VZAVZ6Uq3Dne3KV0F0Dk8v6JP1YOdhXKCJoyM2qjRtGD
1T0QCyXDOBN6jU3/BfKbo8kbYYqIi8UuiiKRAruxhQ9tDJpqSFy0p2M5eeeLrieJ
zhR18CvUqTh6xZBsH8VRHTxL3ICVq8eVhU9vtJWSrHKEuPN2MKJnVEIq1oZMc9sJ
cG66bqYpvB8NUBV4hUUnnDo3mkgiYDBBRj1H885rvCV+6ia8dq9iFW9WPFOmnIv9
NTkkOu2Ku0h5qXOQalhSc+Lzz1iOJgBRzCcw0EobfohLWnPQB34zfI5ssx3iv5nu
c65BTrkh/hDcg9ucfhnZG3baDXPESAB6/bOkWvDYf8y3DGQpflM8bJ1+FmKxyUHL
E5xKSe3+J8PshSoXgSH1JyqXOhvckqhetM/52T38V866FgvkLeTD9irETTuqt/9H
2PW1o4Df6kmdW5X9ncpATUpqJ+fwddwORk6VGLX5Zxfs2VutUhTl9xkg6BWAbOfc
ezLCve8fJjq/l505mo0lhWO85YUhsX+klEGqPe1/1dTBytJNiUJqr0aU25NXA5j6
mQtiGe9lBmKd0EPU1iruEIZ7ft5Q/H+1bkGRJupeMwovg8h4VtWBEXxKLol/6CXI
Lt3X/lWO2U2pLwwvQRRr5Qsbwja6K2WKTT40wISBFho2Zn9Winf7TiG9I8MLn4rN
vuwaPd6jttp0gHcaIXM2V4j6v/OMH8aA3cOHq11Lk3lHCUpD5Dd/f0y133mFlRvr
wBdfFvHpO34PLfy2qx9xaUCCdVtuDgrotUyx52o6ubDFjvmGsUfvrt1pWv0TBcBD
uJ9HngTjToo6SpKRITSpIzQzwNsjeqzhkttYav0aHi7WBUb1ZOaPYPfbHKlQniTp
ca3XqB8XRG9mQUK90vso3GlB+4hXRgkS3miy81L9daLWrqn5Ju/8ykpzVj6Ymc1+
jD0fER2a23hDgVtA7JuDjb7aioTDleQKvcOv3r8uZcamrTiEvunCpbJdzW8wYnyu
n6pzPKcEtOI7LtTej5wVnsSOAYQzN97JrZLxL3KQGyHReYrg5ngJPv4GVS8Xbuq6
143dgulXL+SE3uKxIcU0NE5V5BjOMbULJjgADqUxjBPRn02vAfWfFbPnWWqIPvGO
GbRWVYCx7vTS1VaBOgcA9Smk+lxpc64Quqar8YFU5XnkFe/fzA8cp9UDe71fM6oh
JoHfC93dh24XVsZCMEVrjhroo2jCIqRCzQYz2t79DIFi60JysUtzjpG5uWHnf782
/fai/xKt/D41Bjmj/cUdpKY33lWsPpgne9P5Iw+0yzz+ZG0rPkYflSG0C+7kX3m9
VslET3YfME3bqWX/jitI14Ks/bjtkMYWQXwuddaDYknm2ZDgMcItDMEIlvE29mpa
dndtT9gU+HkdoGVenYLWPhnYweLg/veXh3Fil4+ZLKDfeGUN3tyObJS5Gn6x7F23
Q/G8Z0JB+SgPoM8w0rqzhAL8rITUSAJgOv8brMbk9EFLMsWBbIIFX6o2B1QVYKD0
WRWrhXHe47uF9runOATWH1dK9qHrDbQ6iYyrAinwauj9BMRenQs58g+HssygmEDd
mSsUTR2Nl43Hn6QnB3KB/IMVbrKwMvh/7m/dct/+1op8AD+6n1Kbc496TQ8ExEq5
x0zTZX1ydGeamkMForDjGq/Hw345/JJYmH/cp8jwxcY4eJCTujI0LzYyzGXliPcn
aG8zktQMZ6hRcHw890HMdUKzcLRnAnko5wJs7c2S8CNOYwu1DaeODYDeUTryCjuu
bj2n5w27HbUyw6UXAGMn7QybiNb2vwcRE+3xlwbKKmPkLbUtroqyciWq7XmjAxXw
OH51wlMyd6vK8QpRCrwfyd7X8dXhXBkbquHBTS1IpVpObSxxDb4t2+7c6JdAe/sR
3oL5W5edqmVlRskTYfST5m8xeCpsVvizx3Y0ZrHkw8ty0UWoBZsP82xjfMex0vym
j3oElicLnVxoHFIIki9OA/YpOvVaR3D/V9FCkyOVvGX88KfvzpiPYeZ9DNuPEmsj
BTGT9xrN3Sg1g6j8CFQmQxBEk+6mGNJA0vM2Op7/MbOVQaRKj+8mXOZV+xuXX20V
p+Px4XyAG25C7L6G3pZ2PQu6ZEap2T56l2NAv42nb2lFF1r2JYsijlDlSb4qLQGn
nBMN/sy8QUgR/ytXJ6Uo9bibYKUWdZGj7on4FVPe09aXOUuyHYrVWHutTs5zw5Xn
uh1LtPTW+FhumCOp1bQ55pOCT6Oi1RoFzW2lBsUSgHKf9okKRJEiMQQwMsQpz4sV
CkTZyd958DOg/rzCIK9i192azyivQfLBznURyELCtszwWxyJvhLWev/hzHN6hWyE
iMksZ85mCr0cKFsoTyBPmgtFWF2p6eBSzJ5GO8MI2YVFNAucfs/ZDYtRf4QVHqK1
xRvOw3fy5n+OI4kdwjRQKEFp2JA+bAlku2yKE/V0Im+UXEipJ8atsSIVIIp1iIf6
ckYGJNFV4Mi8r3cGqe/8hfGF3w1zzhvpVrr0TH7a19cyB1mZYRBArbztmvG+6uCt
CjwFhLUmPAbKAgwt8s2cirApCkpAWvIbVHs68zc1grt0E/yv74jpCoLMJ4QgqLfM
ajK0mf9n6fQllfM3Mg37f10hz5gi6Ri76vUdPun+v3LIPsBGsWgRrjtT/0UjwXR5
kYI3pyOdx9M8jieEtDXlPMTHn+o7HOxUcBsAdL0oVVvrrA95XmQ3LqfHCPjyf5WQ
jjPEbD6tAQWgM3Qtj1zrwBIZP0S5OPpBZpvqPxP5QS/G1JmH63HL8/UYm905qesW
7qSYlbTT6NPigB1FuW1aODuldlloEUptSkbmTarl1OT1GDioVdvXl6OXojkP4BEU
Dch7tEHdtnXmmp5wd8H95fmpxbd6+lzzR+jSu5d9Hwt5fQQKmdZnVgOC8ARe/7Cp
0Q2A/Rx3YJblYt2ay1Jn+LZ6T64ZFiZJLarIC+hNwGdLdicVSpleFbjhuhlicAjN
JlILmPs0XO+FVx2kdeRN87WQwIgbZe25LY7FyIHIS/uk/OeCPuvyt5/dHjFA4Why
sjR+i6Ay7iuMHi38/1b259rYGg7Axkt6+M9GR8b6LQxPFj3ep4oRvy9u0FOsAYAy
v2nyijSETe5Hb0ws7SULImbT1Hc5ss6COyOFnKWXCqRfUpXgHU33RJgXJ9lNIn3n
m5jxrO9k5ZxHnLKWD3ME/kFYh+8JeQRdTLHZyzHK9RLArlq/s1TDjBf9BzGRPgGJ
IOT5Ia0ytYFHjODipcTc+Dyt47Ii4B+bNtXSCFNZGl8u6y34XxOXw8CuNjPUEB72
0m7Wu0lJlHkuCzuM/Oxz1L0TsdyMZAZKRrLpm0Glz1ef14imKsE4lZDUBgkYkCRq
HV0/V7moIZKX//UIyhs+48mSJyzFN5c08IOiaL/Ma82Nm3XvPk0/C5UJcKYmPc31
w+BfZKKa6p+ZuJ0zztpjw/PumTL7nZc+kLUPy0lavGM6wV28M5uaucp/c+d0V4kk
4qHSrsI8ltTcK2d3GfWviBjQm3Fsyg5e/J7LvS7qwomoIr/svbx/6BIWdn3OEocz
Iwu6I+aD+Ep0upP4aeEoPMB72dMswKyrZ+7ZHFrC3TCGn3ut3ePm0UkJbeV46Bs6
L/cQ2fZWH4MpO0cNzImgqKodVszLR53m2rO/4S1Udc1na2gjykaWPPtHzHRf3Oke
xDAiwSTgY1sqw62fbqR2R0SlcIxulWUFv4qyOB/ur/7Xv4Kh5bkk4cZzFgbRa30L
MxrCxoH/G2qeP37EkjzDjdvLsvG3vIu1sW9TvSz/inKuhms4Lr3gxW9GTLpDxrcY
BHTRzZ4E/U3WzpPGS7/yMHIy2QpAe1oL84MAnjs1tGKbkZRXWkwU1ev24HXe8BAW
19EHzSMYvB08szKXrAQOoWaYrkRZ0igRv4pix3z1B3eLGpYiGY0NYaIBynqSN9XE
vO7RYjr9nRAEkEg73Plaa+fx3Ysb6yvZbulRkmlCBqqwb4YFfPFDFcP/h+W43/rN
lMr4r9VDz5WK7cPQ0gi50XcJCxuFHzZnVomd7QOXRraSMT6NhyncVMtfiKop2B++
Bmrw1NNLO1tZ1ZwTa1UoW5F+8VEaEax3NGXjAIZtayCbb2B75CV07SlSMQT97bsL
kEnrbUld1FleqR6+M0l4mdSyzqQkgXHIjT9n49ZAVI01WUV/sVB2CxBcjv86lduJ
kAHu3+a/AFf5PMqIhqhtL7DlJtceIT+dRP7USerEhDZbhOeGXZy05MvFqjC+wRxt
SCtr1jYkBJhRLuuY6s8s6Wg4fsoiaiBn/HthZfehIDFVYmVq1XEJLdrECTpMmDWl
Xs9hhA13vGdaYx0twbAwTBEV2CNPOsSHg/udxq8qrJwj3Zxc0wCnGuEvm+elVXKx
Pm94gicewT3bUExlisIOSk8QCpJc6+petdMdq3ZxLEPSAlzZW8qEDRAAV4UUKuzF
UrPqiXBE9AOEKWfBKWVsdO2ot2l6k5urBxHNy1+7WtoSJQs4NMa0+sUeuemiAk3g
FirxD8QmkKoW6qzpqfiaui+rojszMtre/NwIiRn9V5vuQAdNehd8LTPe875JExtC
RjfXwVA1NU0LkzAnPxd+hUP9tbkblf6MC1tfTPI29L1ihn3oPhanliuDQgERQeIs
YmZ8UlgmFvBZ4RSCCVjfTcevSMTYmuyTsJvoeOYfsvMifusdHCO9ubifJisultsE
V2TarNEAytUb5ha56qze+rTg5D6rGBYLEEUpZABBLWAbOCtxe3IaMKzM9CjrR5Ik
2U8OYZPlk+dTKXXwsu5q3YXnD8hL79+XEF+PWqPZxHIdazExV8mVqIgswWxRYZnJ
a2yDvtf3a6oK84goJiLDfKmjE4w3tY8nVmqi9ThUjVKmVspwU1w+FUBWYkWs3jTF
IwYaYBP5yv1f4jtzhQGxMG/1gmHcqkrkceL0RgoCDgmZh12Z6MFNz+AnLsraVJIT
+xvTarJdFKhR6b0rAKUmejE/ODaTVxZv8hIXq2v/0Rxv0qo+MIDbWVMucvP6e5lA
9GvSlve11SG4kqFpfsuh3YniktPE+OOff9cn9GUTGTYu02ppfjTXih0Nnj56Q8AC
+OjN4gK05DwDQeWDKlfxhM/ryniUO3I6HltpUdm1tS914Euun3/weUFlrDXWPhIM
tRmgmW1tLQ0a9xBamAwjkmTPKxuPqzTCaoGs2zz9rvsGZ7YaHB69dCbVWVbA6qac
`protect END_PROTECTED
