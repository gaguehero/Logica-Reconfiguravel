`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
svOqRkvFrBfUvr5Fb1rQOcc4cPZnYmrDxNReDbACMGPY608xJQ4ifGIQYIsIlDMf
lVIfkDAVmnTrCi58yrKEFLBKB+WCQEicsY5PTHOYNSb0UwLriiIXsBhkgYHgW+h3
gaMGllzIz2c4A0kpVXPjhWAtG2S519ItEbdRtCsjn6NPeHcBY8x7KjBHunuXak8P
PB90lsEJ4wJ2zdAFQ/4nLez2K5BkBhd4gQH1TmlzclxljRhMJ3xWdK3iUQPHaaZB
9j1XxQe2NegbSsqJ6d9qY5dzv+fO5bvPfpob4Y6oDMGPtKkKlnZG8QXgHsl2Lngg
0CbitBdz7jPnlxR7kyn4iyLsIyUz+28+JNQjT3JD0OX1OUspVPhhUkiJoaNPd4hJ
qKvHR7Ezbv+YxkEHUd4F2a/2qSjU8T6FCWAn4jFBUhZ8qGYerXYKVM3QCifGhybH
JUT+WwgwCkO2iWJAGjZ37052Wa6KyzO8ieL/3vJ4njFzG/EIWG9YNU3GyXXK1aGO
9HCXkX6JtVXtNVpuHNEXePCAGIL+2EmcID/JH9jM/3wvx01m5fitV45VmIZjg3VC
Sw0toDNYQpukRFxwYWQYWwvZ6KZZmhVxONMLjmFYfFZWa7MZqH+AHZo2nGFyj7jJ
fyT+uCVN5T/ioE4yMqHra4pOlZPxaaGwAWbFz/TVmx9wU60RiIgf3m2HRPyiqUs5
VJ3Xc8jA7tgJKT1amwIGC/QJJ7u4PojD+PpnywK/R2QDlAh2F4Awt8pPaRRBja/c
enBYl0fcym7fwV9MQ2yyiUBYTH11Z3Gn1BCmZ5avOokomyYOpn7CzgmgOPNAhpXZ
rVSU50hwkRxzGs01aA9zTRZUagvtcLQBRlRNXWafEdP3BRadCWOalzRMBKGByuTj
Hy9jRcI6Kw8Ezde4n+ujiHE+jz80P8+hzZdjddCWEmp9H0Ryi2xOHdrUtxe9a6sn
JyOLBa20JoJCYeA7W4518WPvNSWZaWMfoI9I/1ac7uL0zZmrlJRs5D9y7PI2g1Tn
XZyhLTKK4955izuXftiaWoQyd45qwfgwNy2Kqtuob0z3HE+lsU6DBEO/zRDWsVzm
wKqTf+IlK3pmuUTH8YU0gJqPvpR7Oc+S0f6tBieVJI4nHFXXukIOWVVulIe6PdCL
I5Cz/t63VD3obKXOU+EeDAaO9Kc0NtPpCYS1e7nbfFncBt0rDsnDz30YFLRiBswS
e7DYQoLcbkIxelWVOvdAEk+6HIkEnZyKao8huTFeS6D49eAsFI5w7GsICY3jt1U0
6kASQRqffxduJNFPTfjiRbrq+6WYaM3WEjwxTtMSS89IKPSb9JY7jF7oSizz4Kla
bKzY/URiB3RjClT68FoC5gMg0JvVn27ol3uutttG0nKn4rFp+3AkkySG6obluQZq
zXlWYtjR66pQCED536bIgUdy/2hZ5/v9hYldY/aP/XCyOM9KGD3T57vzdk4WFAz1
qroKPvtvzxDIDgpe3yA95DIVoiCdZAkvjp4XSKJjHp9Uo+GakM9cOCJ7dKPXvArx
iQ/rJHLmMpBB9oMg7ATWcjNrNQfa20PVFkZugoL5qba06R3JFVi5zfCmcrM8s+IN
GKr0+z9G5fhbgzwa10G4ojtW+RVv+kNoT3AFpl0+LjwL0nuzp8jJNcuhQvGHKN/Y
hOF7lRznRlb4yuS8Xqc5aUvTqXU0CNSzbIqpt44KTyUboWmL4tDQUGJN2Ph0noix
84jsqiZG5EbxE2qb7aKnk7ZsYyNy0oJlnQJ1SOMOaVxWX8C15Q/Fo7UwKFW+N9im
h05o4Fk64XViwmwHYNvqSxtFVITBF/pXjsb5MVxZUo9sO9Qnqd2vhnQW5Aam+7eF
SS9QsTKHvCzeW22y2ea5A+vQvegueGJc8lNcKu4JCKc8FRwKFb4VrEL2KtKLRORY
AqDQtsfyvwP1N29zKDkPa6ZrhOG0rFXnh55hZygVbkLJrgwr5DXEV4U7jR1hzGBU
1LKGXTtb80j7uy9PkIBraVdaa+mP2H9KsPen1tr33IsGSOjqDY42W6abeQtaMzgc
wWe496CyKRHFicnp6KRS221OaGxAxvIX4MnVR4OtA1ENQXKIxFH1pnfok2Vgv//R
fG+woQzgmq4/65vfouQmwmLvGcLzrd3tppqu8w38B8D1Kjn1BtOIOiZV5un6KNTH
A5coes7mw6Lz9rZCMtDW6KIPohGkWHlzwVMNg+ZojnwExb50diYUw4SJuWPXQqwy
Z/WEhiZhMPQLCx44gU7MqQ==
`protect END_PROTECTED
