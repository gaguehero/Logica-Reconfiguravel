`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1ydTJWaATyQU0yWpzx8qe77voKoIkS/Vfq3kmdr7yxFO9oIN8WPt0g1EyMxO4a4
rX/5Gz6BVa4jkTC3DxUqyvI3skc2PieIIsJhb23gwPkZGDzksKB+kujQLpTZ9zhY
NGxmtKE0rSPJ2P6+MAxtlmHgGYPTMjwc6jCruOSRF/LFeT59Du7lUsCiCGBsnBU+
uZfqUUg4MQp4XAoEGDf9mqv7UzWsDGkqg5U3LST+J7gg7yCeLrNor0MqmYOApMN4
AiK6mCmAJec5G73CxaFVBkGSMapZPYbHlMQBtQ2jOmaRz4xMb2V/wWIvV03/JSDl
elAu2xYx7AX0TVsaGe/GA8mVOAZYzRRNHTPi4nTb6pukEqXErx2xkU5v7oTowsAx
XyDs8+CxTUSn8dL3f+Na2h4jZ3+FNRpuNPufrOfiYQ9TuxszRg+9LDT+ZIR4NGzI
n6TwizXe5ZcfhbL5I4LGxned5T+kuy8HR41ejq/isOnaFO2sZGPnQSQOhbr6WVzQ
EzdAGARrLcJ2oNtLYI/45IDFvsfEQme9ba0twzkSP3jnmTetkrodOMC6XsmflqFR
z1D1FWRYKske3tysQENWMAqMzNrjN6cVySvgv+uHI3nC3UyRcE9Dk09ZUTd3gzU7
E/OAV3RUc2bpqqS4SNfXodFdiXXYq0hg2iB76eDl2iiG7ZynLvbITfC/0KForiS6
iZ32R9VAY6v/2rXRFD56fVPy51YbJSZME3yb52qgAdsEin9ggC2ILy3qONjWbK2p
ZBSUFkzAQgXYTTBMKSAMoVILGKZ4ROxLM7JlMI6QKfd1ebJeuJPFjhb1H+Z3xgw9
/BvNKKI6/MFvfZ1WVpnEzIfucnv/OSKkNgiUll28NVojqrc2GrmOqfsv2L2894Ni
5yNGRxUALPxyK1v7GDcJBNEWauSgntsF2AD5B/HHalTE7A6PCdBpCAZER2b/cR3c
wuAupOzswZReYh0tCFPOi1j89J2JyfNTbAVu8mcFE6PMwQ2MQ9DxZj6/OtnD4BVC
3KYD0GHVDUuKrpc6EH/nGXYwpI49sSqUMfIgTEDu2qKvdZGUyccVb05oo+NZ3AdV
kD1ifFLqHl6RXyUpD2Qk2autJcxuZF5OAGbw/lB4gvlpEUmhehT1VYOIZNTdFFbx
jP0NSxnyEPua/wal0zCprA2p/rXlzF1VbwYzjX+xCVEKjPHC7/Hxk49E+JIC6Iy/
03a758qcWHk1TIR7fJR/1wcXqAnjpufeTNO/PqhfvKRDhZEmvQCgzcUWUwbrnkEo
7EA2aNSmCOwis5mCNFSmSVJ0PAYKsvo/ftGxlgwPaHJyFleaGgxfwZ77w0hJiepq
dTY5D0bEqVspq0H++hxTdBupXaiv3fNk+SagTDl8dKbv2MVGj583A0Bj23CbstYm
MMlFjXfYMBCQMS3GtlbhYLcaxAC7Z6+5MFQOyN91IXgd32NSUGpw8Xc3a7uHK/4W
y5a2TPKtUKwApB4R3Kiw5USa07s1IXQ2z71ab0KQRDCvnZJOvLzKWhIB0HDIWsll
Ha5qpotUImlbkRt19Hy1igg5CkJj5yl4JfIUFK+9hEcj4GcmIuLAnsiQPvKwIy5Z
PdNUvrrniNVyR646tlGfMD41pA8LC+pX/LUD46sQhfg3NmSFE8AE2fmCgH3UgpPL
RoAEyrDpZxkxIcrXGcF0spodoW8a6+ZFabQwMx3RcYcJk6z7ty2r48Xn7zKBc+Pm
JWxpipct8diy07tWtPVZxJpCN6U/vSus3B9ljt83K1xRg4x+jj1AzWsvaxTSfMH2
bfKaVrI7RihbhfHguEhHeomVyrKnIc+v+BotFAzUJed5nFfv2w0T7vXUsQidT2fj
evEsrScWBFwJtp7uHUlJNoytDzDzU1V5DifRHaYvwDUaQRuq/zV0XVfhi4S5XqQE
hgmyzOVAimvK04kZ7zvXxMcGT6oojFSDbMgrWVNMWn+WBcEA1L4SQD2J2/V/5+ar
TOCwmA2dgS6lDIdzz093BPEKUuYG5Jp+eWye/lBSJRGfXZDbcs+KkTc6eDjOfC+7
4xUoSjk5dfGI4eDQ+Yxi9QpPSDGnJ/dVM+0HQ8zvPetX3T5yKajwecgUd7Yo1sXe
OnD85pzJ7dhkZ7DqfnQ+gmYcxxIb3RMqfYzN8cWIQpdENPFDcrWny4kKZwdHtGgr
qcrNNCUoC5A4rAuDT6xIKer9ZAp6M+3nyH1Jhx5Ww2pAVU5MlOfM/l8I31OUZdAd
PeNGldcfsIF3g4I0qhjo9S418eS8xqzPbQQ6kOjlalget8OC9zOh1XiVbWccvgzD
vNnDS9bqRC5XT99r4h/omzBUpjVZ5FqzlDiLmG9IkJrc3n2WkDRmq3dwQXEiV7bz
A7hBRTmv0Wif2cbmN1tQLTItYW/KjCIyxSjvLWpgUU09064288wBHHabniquOmkY
izEIU33q8uqPnJYhpIj78lLPM/9Td8Z5pUR94/nVCz0nv+rjaCcMS6xXTLgsTZL4
6z9HJJ3n5usVBt0pJi4TJQrYauOvCDRoIuxG17cXUTo1EjzdhBSwpVVXnkMM7Erk
9aLcEmOUZOR9FcobZ1f7/4/3JCxoIPmymImx/uj1PFWbaxKQQl+PLPbp3EGvbjhD
LdPr3W4Po4JX5VoHdyYKwSEwGuall1PjZHsgXTwfiybYvgfyXc7yLXpIxS1AI4CQ
BjbNy8Wxen8xcq221GZ4HjfpCYQSQW2lZ/3lDAhBfXHMqQJ01t0rJteXNCLiBHtP
ywG5c+HFojBFEGsoX6AonnOaRjsXF/4ioSZP5NtvuwUGGSFMsc5OoJUariD3akFV
QltAlyosU1JKj3NS99YHvKOiaJmRC+hqrv2jrlRR9WS7onbowXTc/YTGGBcHffIp
4D2Y0x4QfTxCgcmvUjOZmN0Kcem6ZQCXUtuaAB+tfZLMkRE/bDtQaxM81Xg28WJe
cmTlwqYONy65hILMlrPH8ESGLCaBrDOZx7cegnzgJhxvWV/Fpey1qtUxdAu6yVzF
y4ah19Oj2aibDv1g4x7rW2lY/HwAone5zR49hdyW1An5gb6cEHRarlUWICHrcKuV
1mF/prlRPUt7CLBSVlbltT6rx63sjDGnQcXK+/8x10mmoYkQjufS1zkzUFfdZHbC
e4/u6aoltQB+gdfKF6VqjMn2cdlAsk4PY7HSnCzCduRHrha9Z/qljThBe70PsZjl
xtuaQD2+rEsz7B1O81nHW1t7vaeZmFICMHukf6fXQAhTjNm2bh9wterEyHUZ2UEl
2z/6R3N32kMRvXMuEQBvV+XN+k6Ea16TPedDDrWECIx5OOZdz3xpC2+hyg/lLVVs
K3ke0cRtvVSYf05MZfixIkqhuXVqVw4uso10UO8qe8yVUCrT172PjXKA4KGcKfQ6
oOiApl+6zluVaL67pqV0BZYaxR/YawqzLOwfg/xUjH2IZmvsi+8YkSJSM8ZHEtfX
NJtaHQyBBinSw11SprVkQxV1ItIYMFxZ5HbbtPQfgo362uTZ5a8UF/udD47iJd3X
6c3m/JniAFayWqauSeLer/sg2MlTtJzNIrlR10r/7XS33TwLAQwoFwk9J1JRwUyv
4faDVBtVfWrNHYP0LJnr5iQ0JB5vqb2L244oSpsy+vvuimBR2ONVcMijAc+Xy42z
Ol6Jiq5D1wUGbbxv43Xy0hDWbwxyxY7AY71OcGK3TfX+BcBe63Zd0rib75loMCzL
jFtc8aZOQdBiYR+Od/6k5P2LqXHVWqTKLj0X2FnDzVd3krOex2/r0Tpp7glVx8Ej
sWsJKutSvSYUmxgDTmh5DTqcOV80LNfy5QV1FoEStp0SkkWAzutqYdEtWklQjwd8
5m8nDwtZW4IzjsmPXhyFwqd3xp1KKgGqm6+nsDnXB9cvC6Ck8YO4fPN3pCuQaBCj
JAIMpRGYn/qk5oedyecl+eod9Qks9FvT9RJjQkTuLFfSrgnveNuUFYa4Tdj7bbiK
iYd+M13l04mNf3xYD9gJYGSatwhJUE/hvuktTpc0czMwU526WdKzDerALerMCMS/
xWYnrT4YGp6/rbvvEP14x/+ALaTIytxh8b0Uz6PleFQXryokE1yjFu67aZAEHt8G
FyCoKl+RJp+fz8J6758fe7xWoqSgdIyl/fXC0lb/LRee91DwLk6QEcf8HkawFGiz
+Oz4PzZpPcD6czzSjKwOiyErRHJ43tlykfwqd/V7Zc4FwEM9S9C+BFGTvAqrC3zo
a/su3TbdqZxCPKWRi+u6H5S4KEfuOlg+/dSZSrUcCvaPVwlPFkWKiCuGcewp0isb
Bly+kG5lgMGNVrFrOnJRtTtOtEX9ihrwhVdHb4uW8I2EQb98GRfTrKu2iaDuEK6K
YYn2It79gHzdup7vb4NUZaT+fwEFqvLPec87PNLWiAHrqvYtM2navWv/Fb7gBPMf
HmqgWIc8ytpBR4p5w3jqVzparz1yYTdiU7stRiLNPDmQUo4g5BEKZhEVupJy9ElJ
a7lbU6XwsYhe51l14d+/khT2hTLXbn/Vy7DI9zStep5+OuH5L6RHXe5ORohBe4NT
W3009djsN3SDd/J+C844oB+3g5/yUuGpw/QNIOajdd0ddPRranWEjYZLwqToL7ci
IBNbvTKvzTWcYI8TAfkJYWoUu8UOOVnhvy0Pdr5XZ+V3EOvsTq/Bmn6O6plKw/DI
f6Vyp5t/+Kl1OAftwEPR4m/6z3AZ0Z58oeFrEc6PoXApllJ8vn7WAPmrmKOjgA6h
P7H++itV/nZpfaOFA4vYAF/S1whPq1IU2zDw3wWYylbjgHzfe79HMYLeGIqws3cP
xzOvzqaP1N0D9q3hN1Wbl2yAs3oKDx/nrMNS/hhywQzi9yfdMSWeHZ9xmhGq0cPp
YgQohkMXysnLdA10/qfIzS9Q3gHPFgh4RaCfokVXi3lr9SY3iUhwFfYYFG3IMEYO
vgG3Ma6H60DgdaXH8ptXmecoKXQ3VHI0rz/ZTTh2zTBkBz+93eu2aae4rs7RieVb
mZssMDi4znqvsLKxypQHXi3Aw30LSH522WEghQTCnWLABHIzakvD9qa8UjTMD2Mn
4+9/jfsUvPBShnqol1r5b6RGGJHM+l87mz1fT08ATbtXPrbLTISgQmwShX83/GKB
xUcPYvPrfoODE5Q3PWYAHVOLKd1ICpBc0kiftJDavfLCyQhPVtNu9NegEBrYzTbT
pKHUlpPT8YFLVNvGZs4DoBs7/bJWbyArdUKLhpORANKsMiXAPKeGNWnPAv0AZUt/
yT7sKd4aRdn1kAUEbwkdsILo/N/qSBXmU6okQohZkPnYJBjl5pGqNRQeEGVSvOs3
6WvOfvFIMoBWtbmnRJtlp4ggfhlmM2jzXEzRdVVjqAlvTRXjUlo6rDX1xshLNdNC
PXPlsmiiPf/SDOMOoGubXsdq1XIp6QzRvXe2v2JlHVgSEwyAAEuz/PKqDoEUrWlg
1Q3CCl7myOSeOnQ78US+UjKN31RL3RSVGoaZfsao89qO1OtnuBWhflGD6GZKn1GE
3svPFd3ZGx1M2g362knHq0hK1OsoDrDiSd/1+1gftPeTz6LuMPK/y1/gyu+q35ar
Bpd2XX6QT8M/a1a10KEv9NW2IUxprzzfTT7xwyGi4mz4IL2T0YIOtJNn9aQ2NwDz
961zuIh0fUL1vqLB3+299wrFQXVrcKBeAB4mfGX+axiR0sdBAl3remKE04QyY+ow
OhTUr43KUG+NLlyq3VccRVOMVrTu/63KBrUpQg7MaQhN3d6RydHUr2grDQ0TfmEK
JA1X69PK9F01606bl9fcYtUDZlURwjImsyAaXr08irSat3AAEf+8EJByzjKbdSrR
qeWaT6yh8SfWicNrB0lL1K8sulb+DCyIg26dGCrsEaRVv1k2RCMtu+lMOzdx9W3s
06eXON0FyWIdHzkQXkObkj0Dx/WlRVj9zem1g9jtxNvlschS9pjrkns97grs4z5w
NSlrEr+wjJKOdCGe4IA8TroP0VDhpCCmWedRK0IQ5JqOZ/Vq14s3RU+YZG4Xe01A
m0CDjSFQ6a7yqqsawabcGCjcAq5wYxW9xzEWU9hZxYTMIEs6vteCglz0vWOZQTUR
tlZGQ8hR/GoEMpjhnJl/2963d9e8lQ8RgxCsq3d8qWjxjTzDfvM5WCfLkBPE/WME
Lje/fLGOlQTwpE6znv2dWmMRzPPdJEiwSIvO/E3UjgY5fabvoOz01lq3W8GQ/gbd
SnDb/iiJtSW15AXbr0JET82D8/R6dZmpZBgUpzFE8PDASFxBRyS3Eq1krg6dD8C7
9VUcVCYT/Gl4pGntSrQCf6qwuS98ybibp1M7LuSVCbEo6eet1pDFd62u2fkMXf1+
TbijccJLbfXCT2/QckyHAB+O+tM+YRlBmaMjdwOI99fO1bi73+aokpqggd6MIDuR
+6xDoTRUEmUishPhGKB0g3V+XqRGs2sUSQb/Hket9Piy5YlfinwgOYscRyvG9bqW
hryo2uiCIhXYAf+da2iSY7vqVT2wIENMh6u4fbF/xvHhPFRCKBPHDB3psLj5GoeP
WMvoXeTSdUPjH8JZUqkFkGMuFJB2+LFFFrfB+31XBw6LWkTboSn5m8GZHbIjt1mc
yP5ylr6/xkvADFfdW8GgpHjJdiex7ql9jySKc4PVrENjXg8Sf7djCjnHD4CtvdFF
nVe6PQa+p/sW18NH4lJLGD6KZOK0XalmLPylN22rTCKGYuZVn25cTFnJ39YQN0N3
OlZYLZhmnlXFvk9h0L3lsI5gUZs+iEz5tIDlSMtbBE9r93Ybqi1nsFKp0ISXVT4f
YgQayVmiNFDE8dGy/H3p4VCw96MJ7jIo+1SrJVLb77+faap/6zKtdUZxnMHCSTIu
i95CiNfwrQ9KIphVlvB0Wze13+xaKT58fc3nI5Ood2sepEUUkVZZz3vvCmOjtmDd
TBi3YRGGMsuP5O0RyvD4lWIn1mFUM+95XaCSW4hHEux04pTHhZ1FzjqblRagx09l
thaB58Sd/zEteJokJwyUzWp/9Z9KBOuZaOqlKsACtAhmMRHLiHTyr2pbt3K1bnbU
behxy2f7tZyOa7LNx6yuFsDOyjD70/W1cKtk3nl3QwxK6W19NplcMkCFWApkDOX7
8Pyr/D6ZBU4sUcFAbmpFqb+9TdWjVq7vV85XUylShKHp44FMbZ7RrM/nboFcWkU8
TNcr/ARKwhMlZBo8APXejYa2niSuPiR7k0cnfujyGkRU5s0bfrr6P9AcVRXa4Fra
w/QB33Q5yyV58zJdbxNTuhVuBuWJNn0l3ybVAcaher6O4hFSMnX+cZ3v6uTgWqlB
+ZHJLzCXGN3FoqdORwE6q6J5hnyc+NrUSr8NVwqK0vEO+BSQnHI+Xa2Xrwbl7lOZ
R+/pi6by+k/A6IFrbHMkRQvk/IK2i9ShNR/bDrLnyqCXYHYo4GWcuWTeBibesqR6
cz3LSQX75ojR+F8WUbPMAg46Nizr3TaO4JTMY0jSsFSV3VRJCq0+sbLp7t1xxWM1
d+ZuruFQE4sVqfa/mOGOLRevSWzwhsmklKgPqerB+LGr5pkPI6N28lLsvNGy7Zy0
xlr+ESElIzVLMA6mBCSJf4cvtourm3S/DE3i/V/lSyow+PG2Vv+v0honK9fZF4dR
he4Tcrnwnj5WaGXIn5xcBC23QvtOSJ1CQ+ufBLmhrv0mhHu5buix/aPJ81id2Ba1
`protect END_PROTECTED
