`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASIa8WBvA5KXN2xPLkg8EkfJ4IbUR7LY611loapQfXbHBfjNGUJmJ6GM6J5e7pCF
0tGP7tDFUzNiEkOC6FPJajeIr1DPLtkpf8xu8ct9sdUbIKgX7qK8ZEvyJ+mWNBn4
XMYeoKer3OOv61MAxOutaIgJxV35BXXXx7ooVQlWoWecF6rvLfhj3AKF6ckriL5f
ZStQFdIJpKSDj6yS1XJCKPqnaB5S0jLYUnp5V062AJPXeWsJTMS5qBBEFadKjsFP
xvIpXqn34TIf/RGtiE6kDvSOAfNp5MHMUgnZiY96ZN8/ptG1M95tbF0vL4jenbyh
dH/xOSE0WD3/hZCFE1id+BJf/aS8KMCzoVOG6+KD0k0dlue6SQOnNfdxWEVl++MP
xZVpCVzZOLk77izSx4InbAPvTwfOVSAEzodIS/h6FqHFMyJqpnvMagfJ098aPv0d
tHR5JFamP7vuCezpw+VCi3MRU5Ht9IE1dnqPMleSzUsZ31KPZ0e0vyixg96w1fRL
jJkR0QRl2PjyGLrZkPjtYE0WEa8v6mq8ncJu3syE8LeJZDbfZnsdMAbqWiyYm9i3
gGxbOw+ji9ZVwAOSLZ07wFJHoWv0R7IS5bm0fwHABtGLJkgVRZ+N1V/A/k14fS9J
H3r7/yA34O7oYTAyTJG680tv2EpuWxlWQXnB2zOK/k86igCNfs2IKBIz9owynfgX
cHZFqmnAgTPywQx+23cps1cA8+kNMpum1fxFe821oC+qTaiszFwMEavTxfdB8bpt
nlsNjsPp1/T6RCwK83RvM00EWkuS6C2fEn+iD+h5D6FZyyhikoGw+E1bJ6qyHO4r
U20borHyINl7g/KS3/SkIn+bibgDWHoMJXYMiejCEDqMjy7g2MT/Nu+vku3qtb2V
3XeXCyi4en7iTBDDhJXnPVn9MY5Jama1eIM2kEFU3kO5frVu26Ku11L7ZHUVInFb
7dyEr5s8BhLOzVuZAnCMDdiQwGxhYDtOUJusZJgvAw/f+fXo3W0gF/29Dx4/7ALI
aFcpdZRBv86nK/JD2Wk+Yju9rQ/F1bzySq5QrkdS6LwhvIKix2tMp5NiWsNTWQS1
bglUtpEuD+cgsmvvKsX+heAfIrD5GIYcIfxBqRRxOkhn/RdDemz7LDSB/0ltCQSk
xdgCtJL6GZgmAyMhuQhaQU/rEwo7w0UOYdm3NMSV3nOQ16e4oYNyUr2ZwMbsI8c8
/yOeenDkraieolIHlEgyWGep8PiHKcCVZXxFLKjnARI=
`protect END_PROTECTED
