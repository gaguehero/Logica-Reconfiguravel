`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02ceDctxO++smtD00R8jsUrGBohtmkgRQVlA2r/MQKSFys+4UPBfqZ3jJtWKR8Gh
02Yuq/4mxC05xncLYF7dcStEi3FOtb5TMiBpguwG28jhYTtbdgJkYVu0qYTwxDD0
/iPU6+IBrCJjpDnX2kKw9b1PeYR+SSYjybO2YO6Dk3eA10vg2H1yeEjl23SDwX/O
uv/H2gdwRTk0k9TI4CncW/noTymDXr/XGhhGkif1AfcyTzYMznzrP+C9LEbMCuhz
won9KNOR9SuAzgPioK2LHj79sJOyMKdvtFgYG5WBNlhyYLx1AN5GxFMD2DQB8IqX
L5LfVLWFQYZj/QYSmLCrqm31rOmgLlH8mouFxqnU3JbhR5rzidMCuFafa9T4jKGc
yCp1rWUDScelLTcpouUma25Xd234IgKxdqL1dhBlU1PTVYni5bzwjEL5SjDt5v1c
XOwLyuJmBW/o6mmChO4cirvmmrppNSJbffYOIs677CDhEwMmp8KM0j+pUbB0Gbeg
LuGQGZO1lv363Fw4NEHKRU6LTm2fRDvx4zq1jfgPwvUZ8H/oYF4d2u8Qgby0wJ/1
JWeLsqL2SpD5BqCKEv/aQCmljiOkEqOdxbRAUORp15iwD4RIYkYCP+WLZG3Ue9cE
tDHS6jH2WmxBdTwxDwQrl/cOmelByPJxv2q9n0EUv1rtKa0FXiHeJW0MqgZQ6m5Z
xnZSoPaO4DYsOCfu0j9IE1PcwHUWfIZydbnNmb1dq49w283WKr9e5A/nnTjWwHai
f+nq1A5jExN05+xlfewbMrVtLRgGY/4tgTWFtRo91yb6b4hF3HH3nRJfPtKNJRaT
YN1geZSmOzQxt5TUZmjZ15lvBCKPci81Q8uNF4UGq0/0SqGWrS+Iry3+9AWf1T0A
HVN3EkWQcQBvbd1A7oGhv1PHCJV+7hkOSDwQehCaMFsTfhv18NRXljc/IqV5LKZx
6vYXDi6T0rir/rN6UAiOtteJMer7ugy2ZkM56aByvfebnTJm3hZgpbfgPJEFZdHP
df8zA1wa+QBl7Jf5UYDtw1tD1tlEQqgTo2z8qpF3ByyyaxOeZpEEc6Z5zkWGkhz6
nHLdVhWfcQlZw/UNw5BDmcaWXvSjy0F80uuyg5T0x2A8BS7QMEgkPYiNM8jU78bq
DEzZpEtLDZ0MIeSZhL1Lv9Ws1b3LyfpK+3UY2JBsbuyLaVu1r72LQKTtem+HRkzK
47W0V5EEIUT7IsPaSSf54AqyRgSFKxPEPM1GNnL0hiEGSYHdFhA/eOgIIQymu/ZY
YiSApd2jaSDFLrmhPr0NoLocJ+ENALSbHQSWqCvbtGb4HEuQpWtdTAH2VWf8O3MA
nwi90fzSYqtpnjP9VgCuCjW3T6ZMOO4bGQkRAPe7WApbdpZ9x3z0ZIQj1isKyEM8
M69PZuK7r/BAbCKWnKTValAGhwfV8Zgduholgd73yUHu2UmJ+hHFRKUqn2CT9vTD
G2inlzAx4u7/f5MJ+VWe2BE/NiAPoYBGUmSPkKEjcS3ch5OLEKE/+lHm/YFC/XAm
rBwiD0rfMW/0r1kM5aayuosHt6A8MeHaN3Q0izuDyBGWR0sl79jihlhgOjo84OU6
OFtFqKc6hJFVZz5mWJYUFF6ZJC5YRYYkorzcgGxSPUM1K31NF3bHK1qXiYyreXly
zdYVx8r91CbCiaKwtR29AbYoXgKhllDT/33DuS8BCGIU5Iylb36/u0PEhXYPcLIx
z5pC7m4v7mJxrKOMJc4Oq8x45M5UJe/3tFB5x0psWJzvfBf08WhG+esbMG7jFVOw
zg87kuUKJGTfeTeteYzf2offgGMQQ98u8kQd6wBu7rLJzigwa/g1iTb8KSHMTdH5
9vjkOS+pxBz17Wwc3F3ISOQ8o+kkelwHmpyG5voL6r02NzlZsjk9dTK/rt3gCzIV
JaNaUeKAI5bhh8cGfI3pMz8kMa5SgPJT4hktoLTMcTxivB8fR+Hz62mhBbnIjBOn
PZ2eGXcnhqVL/XHUh2enJJg6Gv0ygjLUM6ghbDBjWlUSmIlvDvhjnHHrLQFt4YcE
`protect END_PROTECTED
