`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HKCFwRdJPURM6pOAF7kET4B/2SQd3SVDgC54HMD3bRTqTHqGsbGFAsPCqf8avza/
U6ZNnfK90nzhvmKrT09vRaeuWAMj3Kue+hLtas+d9wsiyUhqXRWsqdP4DiICH+kh
ofVZAlxa7l6nNTbSnCBsMY6PdqdEYDH++RLdNHZQpR3BicQP/At+KN5/f4UYifSZ
DllwNtCJ43dooK+R9udOCn6QgDCAiDpdz5ykU4KA+NmC2E8utD71HyCo5cHktQfI
Y9fthXOFfG+Jy2oQO2Knm/aaCcuP/Iz8A9QXU3iBX/DhARDT8zeIMSLnfq70So1V
v0R8HgXBlQ4Buneq/IxGLYQ1cMEwYVhKxWsuBmYxgC6QGDRqthq9QZog/ZR9xLe4
MgyaXBNky4VGQ+Gxkchr3NmhksdQGsjOlgx817OAiJdu+jzgmlH5wVVm0RnrdJMh
Qcpm0SJgUf9BbQiuJjQrc4S2Slju6pLd5vhvFiVfY2eGXudN9zUIr6kDBENKsJ0g
uXxABbjD/bv0dRTae/uhzAo148j+lLU3RuB2NraVM7qXnuFqD4u+LK0jUCxJjIsN
lZg2UfFRgEALEciuRjCQSnC6ye0pHg+jikmt9+9F0vfwxtT/XZiVZBc24DAMOrEO
rGcP/HXo5xv169HoTNUvXpBaT2KmNVBIMhuREMrxDww8l0wHQRz6M+7C6FSFuTmE
ZxHAs4QBLyZRCIFqh2sd9tM4ljSgvAmhWAoe6HF4HfJ2OHPukJj2BOvA4rj9a5F6
vssXgKphSH2ajv2zuh+FxI6zhV4FEAaa/ZZu2lBmyNPybjLpRBF5zz22y0EhE14g
SBItxiAI8IffAFbhc2RDED/EpbFaBkRrMfsgsbRw2SDmDfS0lwDwGiCTuMm7s0iW
Dkokt8sBMRkkt+mz2JwnWCSX6EzeTMaah/YfJ5AIbIDsOXbPNRQPcffV8bt6BEBo
pUoAXv9LG+UGzMHv23WyuziVlxAohJqugMhVRL/1VjquEz2qbtDnA+BVO9ayl0wJ
ll+AS5zA8kV2l5RiZVGV22ZPqZPO0du1qq+n6d/1vMfIZEfe5KQUoZNvXkDcOIGz
x3SidFqdRw8iXx1/krtBNfLDYQNR7u/alvBQKBcEiO9TQbVZ87IYLsJuhucSa+a2
qe3Bl8LFqz8WmgY1D+aAtnHBqiA1C6Trr9t2Krg+QH8CXnpYsgLSsGaHLEkt71ES
wIFm6oG3HWMLmP96A/Ybs5sA+Pa9Gzp8KQ+DUygUfAyhYNECJT7snsWgfB4zfzcE
YJpOhnyEvaN776onHaNxyF2RRHpipDkicTNGXDtnjj4smHFPSSgVc+V1RZxrvJ6H
QW/WKa4T+XzgQI0BSPNQOTLZgVtY0u927UaASsEIyHo2Bat0OQx1XBft5DlM2A5Z
W0m4ZmP8luQx4R7BTgpyEMMjCnyvFpFFEk+Aq3oVQAB06s6AYEeaMXVVqUAQm53O
AaEQkXF/XXQRNdrt9uc9VypnN0OvDU3ertCgDMIeemRSkuR9Vglbi1I+yo9Fdg68
yKE1ukqVR6TfmWaZRPcmYMRVO9QBgKiYWsZCCvyJdla4IrrcgF4VKQuJ7ah2uN0F
LRZgZ89h3cxrfRU4bVlm9RsJUQqp1Kz2M/01ikJffbhUyFW94zgbR9hSiFwgi1m3
19chSJ2oLH0Jq7pKVWQRyIw27L8ifpYp+0Z0hd+uwihq698pdo6SeK+PLgPxrXs6
YBpfP5eTSXi6mVAacCVBDljNHXvFs5tfbhntIOMR51fy+gUALxii3hrznGY025ep
K/7ochyMhVdzC/UWpu6A/YhxHo7/HW6RQ6f5aVjWw/nLLw7NacL5QY8J52W7BDeq
B7gVlPOcEJ3On+NQXwwlhSn3FZHiJP3tHoeR6eUUCZOS3STqWycvKII17CVBKE1N
nKggMONi/pygPbZPHTKNtXXyYP1WkdKEVfOEoitiJ06sEJVT4zftSIWr3ogQ2c9u
7pEsy26BH7EQOFK9b0YJqzO1++ide9XJAoQlkEvftEPg4EgsOBZdvvAbuSQSwlg/
`protect END_PROTECTED
