`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xx5LWljen+yFK3kAhvbGZDHWx51/FNCve7UBqEk5b2cqwL/41knvJmEv3HIn0iC
mdDcjy2ku+5N1chsyTJn6BczTNgQpFi0Qda/Lyjoh5SrbrZeWe5+DMgqNVcpKsI6
Wrf+SPaP1qi8V1WMHhD1wKuQi5CESx800+hnoJVmgTycM/Kb5Fj+SizzZ5/huqVd
n9Fdh1IVxnjNTlYU/LD0uZypgVzQbCqhUH2I+tj1ZEdE40bsxN7sHOtfyASvEtpv
4dMm+zeX/vzfIADQ5IlsTO06OJYoqPoDNn+pJOM7dTwL1yBJkcggkeBDqfHVzRhp
bS8YLDS4T6Xz7Q2jLu7irxpyVSQklQo8GBVe2nhNfhtOGmPv14SPg1l0hzCfdBBs
O2fQ4HiLwWoNQ2+BfdAdjbzOsRIfsOgLGZDHleWqLPUnrpklnxo7r6lpscZLPLm7
ULvz9tV4BNDWx87wehUDghZUHgkhXLQQhZdQGrDZdeTbm08h4HM70M0lO2bRRddP
3BEimMA/pOBgxsoE9eLtXqA18BSMZPnD0AiYAtHf9Cv3FIMyZZ3tGG5BS80JX9We
59jhMZKliCLxNLI4XtYzWVsKcTkIBMhfIVx8IxygOqXFaO45EcAzKVbaICcy/DMH
VNEFN6dRxMc3r4TAXggaO+rsMR5DTl1UDV05/OD2nUi0PD5XCnzY4Y3y/sVL3Oww
n/MAJwKqwt41WcwZPY+5B4wrW3GZQsBMrq3FIeKsN4j7HtRD6MxYSCRSJwaz4BSF
5JJ0GW1ajr+0okPAdbJsh91k2wcied+c25UXyTsHnGokoU4xp7CPzY2W8uVWuZb4
jS5RuF0rShjbS0n9QaKs8mWhL09iI5x6CF3m2zcFCs5bjtg4H9neG7bL++SFhZlO
wGFM8EA6ar4D/R4ybXLLfQHjzTaZapOEg5tK89z0VakD4s5kA0B8N7PZoPNlG6A5
MrQ4FlDoHNW2u8N1UrfeagkWFcSIM9iR5xFec/eUQhq9yCpPDzc9QMn1DEyMwdDK
e/8gtQjNEtFleiSCwialO6fQMiaMExc3opQr33nM5SMn9BBKwJiCNd9+WQ2wxEx4
PQbauJ3TWsHS4lD14fkQIAAqxk1laoUfekYuWoAs3pcTTMVhQla6X6yy1vvA1UiT
STPZWD3EgTuHYSRfHlAKDgU//8+aAMKqg3HkqGr9iPRERsv51apwBugXKiQnkkVf
heqB0T/B09o6kGjD7RFrcgPLYhnAF4srA+qdDlwW13wV1lUTA1H1kBfu1/REgDBq
i3/lIwtOkvGdxdarnwSARD9BdcqFj5QYMGJNg7b8eZAojnknL9JWS7gq+MlBKc9w
ZAoqQD03qW83p0TwUXA+6GYoxLFvc/DOwRqlapgPZzwxgpJfVWwSaLLVprYGQ6S8
bZLFsCs5E2y8CV9W8OI1Izw8ilpliKnaP+f7zktOYsiCeVeDKoeF8HscJY+ogtp0
nURZXkz+TELcFwYOycME1gBRSI3yLU5bJhxQwtVHxCw/ZbNszDq5/95v7csBWkmb
M+7uCA6MUDJQLYQNcnjXp4GYdncvl9D5ywgS8wYc1pQu+TbSM56o5W30z04k8J5s
OhjJzbYyXSS8tu/5shy/BUhQjvVQibI0c6G7/UtatRNzJdi29XtinzkCpkdher83
Wr70rW1YVPXNZ6z44NVej6s3yODjguxlmLdgn+bm9I8Qidv5DhThJbag8wTvOQxC
l4dmqh9AMb77bn8yLLa3sJfpAJhOde4HG3w2ciJAjvmV5LERFoAnYIXK7qimKWL3
AG4IUGqQR7bFsGjHPgW3Vw2SWY7AKgSL+dZQwoe8copws4mFEry+sNdZ2dbYlC6c
MSBzP0q5d/oEN7qnRRebvJMSQ6244KjEdUofrBNiyLmQ7o9bMmjCTlv30XqCLXYd
2wAsB9EEIrIed1EB5U9MfuIfKhFNUKgfYYJsowEq5KbqewGLsL7UPzGedxqG9nPy
1peWRPfhC6fNu58cnDjKotlpGItsNi4FcF5bAmVXt7arLMGOwHAJyuvS0p7PfQUE
J8nXelkwymR6ckQdUwjWTZEkBeOwQ7cbFK1K3dCF7l6MkrPt1cu5hrUyNGd0d6cQ
6b6s4Z0/xdqyd9pnTbn0LPaEv4bEzlsVJCZ86td2lpLyeztFVhxJX2Nnh02np8I6
JOFf7+Nk4p5SZmE17m83cuVOmAjs/EkLIcO3YoTEMADnUYihbq/kNPeHFcBl186m
AVI4v5L5DYEI6lIBYcKo6W0qwh1iYc/miNKDh39vD7b5tOLD9C6rmSdAodJjefMg
cG2PnViLqtdQvS5VOooH8nA89r81/XvSJXI6lwcZm/U1AVVPP4o+g85bGzqrn4tx
c3PhqKRlVmLiFiRv/ibjdq52aK2hIG/hKE6z5C2GAUTGVX1To5vw6wBxuWHB0VDx
sEel2XJYEJ6tS54IgVIYvPmit/gTPQgnU/Wlw+y29S/vGmbvJHAsLcr2UR0mtkS2
b7zl/FPHnbBizokvyKBy7lQS5BJ1zlsF2devD/qIi6U8TVbkF2CqKfM1+p2fQiUx
eE4Q0lAMII/2UPZbJLFaPZdueGzTkhpZzqVTPLIsnf79QZ7DMxk7WB3X6kBqbEqK
VNwXLzhatQk62QTBf2jUed7tB2L3440YjuQXMIOX+58926rTi/UUFPm4lSMuc2UC
7Kn5SqdQIa8bnjKb9ReXt89o5HCuqJZog3OLAfKus0mD4p4XHl5OlO5/gejfaeOE
20PJihnVgOaFqy/wMf83dB87WWI1xhPvEmruUiebZmBYjQHfjEyj+Ss1Q0zf5biy
S5IIoNBaVG1DtTedYh1h7ALz6rd9827ECs0ZUzgoUXdt/pKspyFdNvSu+85uhBze
8qPJOUjY/PZ0EeMdiREqsmPC+98Vjy2dezb4PNBGf6G3LFRWF/48bs567vv2Gtzt
1aIjlOMLwZ+ON/j3Zx7XcynEZim8PpsTxbMKCCtpYz94FYZiz/m1puE5+jZq40OR
cwYEEYjPBBxyfoP38OeSepyY7fMi+gSgbaENpeSjMLPdbLENeCPI2aIiRjFJHJF3
XrrSkVNOFDZ4i3jMhUVgATambFr1Z65L8m8HQwIJwb8GHqsLzeSWeqeFWFs9xJJC
B5c18pK+X9/IYNXzv1SeVZ/tSgNFwls/vzAliNDDgynHr5hcdPXbeATJrYfK5u3a
3/e7tfe+GwpMhL/YkZTz9FPmRjGdOT5zms+yf6V6UVW8orDgBkK6i0XLnJAiHsdm
a6Gz1vL4IfBSfYVtEouM58ZhFqDU4RE62OUnTTp05SGaSlk1LcTyd8nvK7980Z9I
DSNxt0E0hz9vRlQo5nS1H4cF5KCDNnunvc8VcNA81xLumvVrFc+b+oh0bCenGFaS
9H5bDwKuKfE16QL6I5/Pi20SbRPbKTAOippaZBwMZ+0QBROm9daiPQaYPTRgkYnO
pk3DT4uMZEWlFltuVH3qTKwMqgqFvjgu30+KaGMoAzyJEd8CWuLWp/gMzomI/Ua5
FjJ+CQcRLH9Uuscd1aQh4St7YhwJQXatKyIr5qivlsWBvN2wEHIIejLPURSxsNHC
fYWdOdfXCPLhwK5z21ZR8v1U6KU20VBZJbrvKoyMmKS7ovmWQPUg9LCJ1cOAj6Xi
N68HGZWBsjlJenp+eWzvwFalnp1luDEhccxlZTQWRWHzpRqESZud5EQwybUYC1Em
8/9IYVXLAqX7KZ9Y4fvya2/bNLeQuUhxd5UyDWaoegIrZPz0ZPsx35TEFzjkiubz
EFKMWQRiYuqo7GPkcNTqLT7p3B6y/y8dUC2qxFF8VI2ct1RXCvIW63zdJh+/yqq4
WZUy29BD/pOHEVQBs1+y/8OchkeeheY5aDxPMRhGdTuRtfbOX7wjAlRA5peFoRtw
Y46pDGRVFNlQjaXWHHHp08CUIFtQE0avhPpR5yIeSGHGoS2C+ctENexV0iJK/Ww4
ZqFpjooqaRtoHqAbdZ9x2RRPfhJlSFNA4cG/JoQm6gCqstjbdWLpi/BXocl0nz07
glt2dtq8fBFsUpiX0yT7y5kVQ7BhRwnmpJ6bQGD0YlyHnkMMeYep7y4r+kZVWOHL
uJuz1RGzmozxfIQ0odVK4zcBedJ+lxwMO2URzitaqHyeO4xRjzbrBevRwTqGF+Ms
Dqcdjwpwy178qN5Ktc27gbvYUAXfogYLUw1/AYCoeO7OHP6HhRlBhu0VfvNlAJ9A
R/7j0ZSXjpuzPSanPq/Puhz1ZqGnMdZoUBqawlGAASysxbosZCa7o2UIUqvFWFoH
OP3f5vIlYdYuk5uFxyefoJzO81ywbs6B1zOh7UKVPRDdhxiY+EpybM3ZewMw5ahD
GDOFtnWM6uFAqmwj5vzcEgTHyPokc0GKomGymbJA772xCn3CDRhhaf3zm4gLw97B
FNOW5Ceo4QaaGi7YuV93j+I1xVsYZE0eI8sBHQBvRUasDE+LgKCF4p0XCWDrwta8
hNBGjK4rMhq8f6NAzhCMaR3Y4I5d/wUoJ1tWTQS5EPpKbttl4gqUvNKWbEAACkQQ
PeicPasUDw8gFyqPh85oAzVq+ZHREcnKMFB8+k9vN66njQdGrWUUIJcwBF7XIRKM
4sr+u9waIoOBTkA1CEcH0cp4h8EQ9mVtRZ2gcBv9bwI4AVkuSQ3I2UzdNahIN3fE
x9Fx6GhRyMPbKon2qZSnHhqEia7De+yae45BUDyvOOATXkLrio8q2i9VYFzznrxS
ij0b/dso/WcKpjV4kYkWBbqncz2PeI7ANezbbs6iN66qzJBrSH2+J9PCfia4i5oH
uw2M5ZHnBT6OCTVed4G3qKLtAf5unTYqz2anNNVjq965XfBg9dutHF+T94O77Lo4
BUi0j69rRy7UmfmbQoQSiRHMi7+J3ax4MONTeyF7EIOIqtK0E6GcTWXM1QgBhK93
sUv4KPqdVSdlwCNcFDmBRD6fxJDwuSla4KGXW+Pxb+cvqcqv6TvPg+5SBQLap9tg
YPSXmud3hCKq0hAlz1YTEg9KZiioJEfn2enca0iCmujZ8faw0i3g7z0vsiZQCoi+
DpAoji8o6pSrr+i9XDqFiojcsxL6rQ7giANZ3RgzBHIuKRINY5EaGBlfDXlXVpEQ
ruY4seyYgWI0yPlVxTx/rBYh280woVKLcTuPmS1G3Ue5JjlSuLhPhhBZIRWhJDh9
Xk2u1ABpKzH0yj6ASIV0mGb0cNasqvc9XZy+oSkvbuqwezX7js9DMvP4UYOKO/PC
Azn7U4rBMmsE9I2Z4QTTVH3fINhEusTA9+IgDASJXwhuN/HLRLaY8Kol3lKdyeC9
2SejfONm3ePHQZ7pPbmT/9BIWaJhCtV3Pf+RlvBL3zeoE8Y8DJB6HEEDu3AySAYV
r5lh/16nY36fsHvRdnxjy5I+bWKY2ZARC+jaLBmJu0V5589lW6uw2hOJvi5x5460
iLJhNPfmZb30ACY5xjvtP4Qcm/F1NkOQaPT4Pp3bTEoveXyJ2uA4Qy/7f2hlRe+k
gDfyQ5zIbXDFBXOowfp1Fw==
`protect END_PROTECTED
