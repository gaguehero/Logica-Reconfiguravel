`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5QYIytRcWtdKelE1Olz3wN8iNIb/IwfpAbKi79rgaJb8iWHzO9QQNnW0edaU3oCK
tYCEaVBwYYbYO5APpG7cxOLM1zUWP6sUUec9oDUH7cYg9mpOQs4rOppxTVUsF4ZG
/cS1bhxihDAjSVEpjHeY3kjGhmykcI9Nd5lOIIJBxST1A02iSL5MplGAYomcIYIY
ZBEJ6Xw7PZTKlkUGKvIcv5CMqy4J5ldvks+q6BizbbAA4JZjGBz8s9T5MYMmFFg0
ak2txnFgyDDcx6E6FijItLiI/vzGu/Xg214cWp37Xki905q0FHLsBEG/FEEc3dVL
CYQ6tohFHmD43UUYboxj2yjKziTU9KEvBVzNddlWJ8XsymqJrFuaT4S3s9GLlVks
oxyKlmQOXN3KrNnnda6G0Zw4KhNr1uEoO4Tx6YP4rUklBtO8U5Q6l0LyvYtclFIH
rLndl9xIGjjN+n7YMYu5+PXtJdYFi2ViFm3sIefzSnC0J1OWbdLQZi0FW9s5AEM0
HGVfVyN3nI3Cx0O5pwg9IKKWPxeRLYmu6zYNCjtiaPoAj27i75Ij8griSE8udsEd
xzOqnGweqiIJU8A4WGECSpE0lzvzNGbDyfahvgLDQql9AZZvnKd7FZss3BQc48Nd
b+wPZzJyPIeyvKyDk/EnfKxyxRWSKQOZVmusRlvcffiOasj+spKrutf08xoUhex5
SAynPUOB9AnzyEmk30KJlgDVNHOkCsclv0gKBYrDUKsGbBAbCyyGhnHVqQz4NpGH
l2SyWqqYE5f75OJ0Hss//O6qLbae4Kl8DcTyT4yQIswzBVzGHsnjTokYfbCsMRn/
cAoyaNgzY7tduMbfViOGcWTmVPM5zPtH6djC02RJCXreNvhoz5KfJFUnpyRwrxfo
soVVaqVcOefLAYDTftu5sU9u17k4T0cjMvoCspr6vVmoLQKy/ct+avafkOoxUQeb
yX2ui1iCInN6knSnhjZHPZwRGQDHYU8EzWAZCt/SKoJ3ZBOFulHHrbAFsWXF6Yye
1e8fecgnGX9AmfFR/UvnCuWUyABah7GhTSFiA3aUT6oM8dE+gfXl4K4n4V7pMYuT
fUIdZiV1qargYCLr5Biyz+lKF8UOMznsmCrDUyPy3vMaVtTM99Haaa4o5wQsCb3h
22cYg+2V6TsP2CTB/WDvqiCBhYuiYUu2sVnIVGk/IWOgYgToPUeUsCS3wBRUa77/
0Lq6jC//WICDIPAIfGQsfWTK/zQ3z4s+BCqN46phyYaBY06uB2EaVtbhBLVzaoro
tsE18Gg+HUBib+pWTDXvQ/PTQsHykkhKUlLTXlXt2UeePCoQ7AwWLuGuCHnSJOY1
7aeeeB83zGQ//6qOjWaVt3J8mZfJ06z2TAZEyVl4fC1o7HCC+zxPLYWxc3aqBRUt
thwFhjqoUNkZSc704y/6wqqGztyFhvJI8LBls3PeYOmOVYpKVvrtRfGOy1kYLJCh
T8k9ctdAQtTABea1McQ7NdC1P8MAg5M6S1/UmdyTeZT4G3jb/TIDftmsTz/hvEst
3DrM9gb1RfjKRmFvsWE/RK2Jqo0lZgpOEvymDBsIvoDjeTj3XNcpTJUC1e5e25fe
O0jgNC1ue7zx7F55smXiE21ytc0wqLYhRyDzdqKv3xe1iO9UmP6wmw7t8qhta2LF
RwZS/EkD6J0kxwrKFyBVeSiwSbpoH/MSABiEnCtEDwEnVidcInFN36aOxr6rgukx
TPCkqEP+fn+6J+deTDekp7WLlOR7AWn/3pxztxV0ANOuyXoiiJAAsIDtmlI/2G6V
PgMAT4KvhseeeBgobQWnNaeeo2xDJHn9mkIyrO6sKxPJMF6VWy/SxF36WtG/rsiR
Od6qc8LqHjKCoW0XS+Frmep4zezKc5k88+qGP7Gos2phTrwfbbkg7ZfrK9+Caaz7
Db57KIxcCilDu6HUhKN3ejXZ/XRSFLs48fZzrQms8Dc2m1lB5OXYToxXT0PDRSX5
gxSD5+smYrQp8oQ3V6i3dph3YrpCbPN885hTtivJ6xHRK+0Ff1WGmTYQAf/43ekP
`protect END_PROTECTED
