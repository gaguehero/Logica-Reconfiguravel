`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHFrPFTzA0yugemQzhwfOuCI4+c5n3IFEb3D7p7oGgFWIb9yMObFqeD1xokn3i2F
WeGFKpDVR/gbAYKXdTlnejrwV+pgo0hsHiIlXXZP20BORO1BmK45KZF7rLWeUbH8
o9c7ck6Y2CK1Vj/NOddFNEFuOCJJHyzZLrNIuag1skg9Lkm0ICVAIwgWMYxbf/zM
WMTLGb4AQA9ZB1ogEiPFdQnUZ39fKfAcMc6jDjXzB8wL95ibnio5bI50yoXeQhjw
uprMTyU/ccDktyZYGccSoXTjow8p9X6lQIrDFQ+YYo8hJhwKh5ClJdgLAnZMHwMg
47zK0lPyusLVpinLfco8xDNDPUcxSqVuF8mXcc5P0I9XKJgfOTNmBSFlpRFUQZ78
dkl/FCe3KlWFEAWSe1jlfp4vcaOnnc7wGicpxH8Zu/9ToDONr6E/Rpus9LTR6UW2
5VcgnjezAac752wzCHDULgSKEMV+igy7U/8nOXE6h6jIXXpHCZp0sUjf8TcF0JXW
NrW+BK2cviJQkOvSVb9fgIn5QA18r+MIiR1hzw93xf9JaNE+vS3DM1qO28oZdovE
/kJ1lzD6BCq/IjXavA6bK6wjzLjg0gavnW4wBnhOKyjiJf6XaAxFqOHsBWSAFwUq
nnJVz5kiavJ/miHPtRXjoYdiqH1G7kaqQRdPgx6QJqpJNBVgVoktdKxmt588El/N
PF61ToPCtSB+Ux6D1lWOZi6aOoOl8T+iPofllrCPm4rq+OQtJ2wggefwVPE/Gv4T
vAZmIFm95pSY9L1gFoA4NkoX26hVzQNXy6RVV5lf3tVGB2KV1jaegPOx6YSAnsf+
wl8XXMRVS7iRQ2tTX/J/CYRKd4tBzGzKAekrbx80fYagEuqKHw8+PpI0HzCx1FwO
a6VnRD3aHryySE3g9rP///u9q78LrJ3JeCwNof5PZHusq7coqcGhVbjjRnVNak26
Cy486XBhj8dikUtJ+lQkpWzpbXpZUoBKJuXV8HQ0KAPtuREbrx41CVHjcl++yxGB
pSou+A+EyKAjVm6G1Z1HWT/u9e/HNE7cv1+GmqOLW77FyDp0iL+l5EGvw5WRs+Ul
qikUPaF7jad0OuOVa/it+tP00EOhzOCYsR2L2LRbZKh7r8XqCQQZTn6poFHmL+EV
HZdpYF1Ejx2M0uUKDSoLjllYI18sp5dqmrjiIyXf7ezOKL+ViPdvCYKd4LwwcLOA
w6CqylsjG74LHeHNAUOYSdQqAzaUrWQsoD0iZ1473HYUZ6ruOqP/zFb8pCQGhIUG
h45F9Rvqi8DUHhbcArWm0oIQ6egVq4SmJedwjuzDW9n9W9mNmWLgWGi1NtFCD37s
2FzBWL7eG5dEUlaHcT99OCadki5sjGLHlL86TxlJgImG+lNlWc/nWyB/BgtlT7xe
3NSy78t2xLK5scRu1tO5slZ14TOQotn3UE386wDbHcbgJAXIK6Q6SNgGIdWwbsW2
ATyT45iQCXubmIHDPeaIpeHLD21INiRPehucSAXQkVpT7J52hDpt4SmX7m7Hb4lV
Qagdp7XP0XrXPwTJKxlN0g1/6zSdCJbc6kEcqaGYvMTNBDkLpSwZogURbfzZHR1k
PoPuUKpOyLDe2esfxYj4gVhdfYSg29CFxa1Nw7GNAjW0FWWOqOzjDjQX9ssgh9VT
iAKt3A3DMOJuZiaYsqj9DwVyly7SFYUmkVuyv4LIp48IFL8oZpHsDTi7/2hHHXjS
wxxUEMf7M+w9ZB/nAHc1g5bpT32hZmxK3+hczgRW8xF4fIPfCGKYCTJe3E0vcDO1
D0xFSiRocgwhlUl74UhY9cf8/fgSm7bMqqtPdOmA53E5mnJQeEzx4KHCB5Lk01WF
ccSLCXt2Gy7SrcP924B7O9xpHROU6sTnjygVgRpNw220wIvw1W3ieCzDULicMNPv
zhL+TkEY+9vB3c1+LT1jTTEt/apznvObWd2VNpU+qQ8GhEoajsiIyoUfjq9g2AVv
5h1MVR0Iky+GPX4FHClN/WFs0t4otWi1fc0sTpBQ7dTg9efCNXCgMJl5epJzwqB9
dhjvoGMm0eVP4oaupcb3NJQuieZJ2DYddQ1Q4BJir9RMlQfSJ5Ro0ibOZVSpUyUg
m52HGsLSVC5Szjd8sW18ovT/Cvldo3LHhqIYOPKRHi6lQwWyQzotkFaftw8/jd3F
bkb5MYaofnHhARy5i0uWGHA+jE8xomxDB7EN0H8upLrXKRP5m/8WWVjSOYmY/emi
iPOuUmDYb7XhOZJ41pZ4v60OlGBbtuqNt7F/Rr4NDQd3Nn6SIEssfMVAtrNai1hc
IYB27nIFW5ogU/3XI+A26mLtxsCjx1VWiT1UL5dOHnKDvlbbEretJszwV0A9AQyJ
QSf5RZE5uqCUT71Ch/7i36U70BQyev5CR4TqfQE8k20TjA+suusLqFt1k+d83s4x
cn+5VsGC0pjlVqpvdPklQ6/I57ey5TwrU8eIeT+MaXr/Iz9gqgl+PwT8UgjoGWlw
KGvaqWtEx7WdhEGUQVyenoTaMN/8g9XcBhkHyZ/6HMMsNP/uQVU7CY0W7xqboXPa
Cvy0+19TcbWETNhQ0qli0w5CO9Ltguqr45G6ep3eJ5KEoQGYcE9Vw4hpcyTzgZIw
aTl476VVsEQ122Jmg4VECpXTw0RnSIbagegjIddGA1Cy/oCstAGZgOGpNBawvbLC
vMdMQWCT+smqbiGj9bZqcEE8Y9FjJYvtT1VwKJa8v7DKxIHZIsULwZmDmNkqUIm3
cwVZlLW5DainN4yy8mOYi1uBY/wQN1JsFeyss/VnhoktnoDwYJP/4ZtBnxOku8KX
e7ocoM+zVw9NVhfHmCBeYaJelCZ7q3AWEe/KoSiFzCpckkQviavw4k+asy7aK6cf
iStflOU1PjpZxUgbTQpXNGpCvkmD1UV+v71YHii8FK/x3+DKJ1sBZXWrIgdVR8FJ
pNh5Uhh9lHXzzlfv/dxiNl9OfoiCPYa5U7cMxjJR4H1oR6Hwt/Clf7whmHkTaayG
F4PY7LLvvoSUc2ATGURZp7by8RN3FjgAO2DqyG3elx575THCdFFnm+BMRd9DcaW4
K5Dpzg2BDayXdJB1F18yEWT0uWxsfiIG1QUjW884eAe9Ok9WW57uwAU2k1sz5IfA
nPsVWumO2TFdO+PhoYXz6RkoW8HgxSEzCKtw9expZ4/y/3dc9YF7SVEyN1KyD/6l
I0cXWcqBuZeypJ6MnA6sj9Cq8m+B3bYjZK9btWYlnF58JofiukEtDO3T57fcNtuQ
doxpB0hOUqi45Su6HEQdGpbl3qS6zNCeHB0EZ5Z4vST633pYS2p54m2sRTWa3Ewf
fgq0jmTw7o1PprrFyKCR9MtKYAokzfXZSQ/Zrx/+FWo/bUnvNCds4vm5ngJwB+5s
62h5APoOrfaoEk6zpIAdPfUFhs3IJCB1MOgBMGlIiJ4vDIXPHcB62lH5F6pHlVzU
grkUgkrZ9oPbB4OFTNJG24hOxgZg9fHlG5OvHHPLFD30UyBQ4CojGKaPKfqsiazp
xEh3L5GWCUqG3kaWlPvfCjBUqLxDpIz/D2YmD4T9raA7lrVgpd3ny0DJ+u0+Z3SP
1lkXdOFc1Bz2LzMYdZPzkLVOgsThs8ClfxCy39k50QGfTjxfrjh6N9oGstlgoxrt
wycDbxgO0I80e6rK7ecpecawvjuDafOBJxhfV8TCq0K9N4V1QJVV78K7qzaF40k2
Hl68QcRZs9he5VN2qSrNL3UwaQvccxRiugD2u2g6J4xVX7gGRi/kii/os8TnJHOu
uw8cn95vHqZyB/uHpmxv7/GK9iodRqB3jMXwDol5iz++MEtEuhSSZSfQpXPRSuKg
ZSBdDm+SA/xSrTdkmKrmwwzsY0j0YZKw4AndB5Z30IDcOeeoHyWBLorlCWlao4kZ
xzOrlCovFJBYNWGfgoaqaTG27v9sb5H/caXR2/ji8aNtlfg/em6gUk5v1SZ46M28
4MMzfzb0XZZUuF/haidWwTyBYYbg+3uhHSVf3CIzJ1qyH+M5PgF3D3GQ8KtkmY16
Pb1cMg1uFyLMtAyanBApV3B0IaVfdQ4OpAGQWNNR+A0V6Uqoliob8T39tkpH9NIK
S2Sd5hqIW+Bs4/OqXN3zRo8eIDSsQFg7lguMjJmdiIulxPVA/giZBHwY1CR41Xzm
NLuUYuJQ9YrxPhV075bE7pFWTZIt7Y32rBqjT5SmakGeZ68Q3z9Ki0KLxfbGkQOV
sDFOFI5DuBEdMeaTniJfR0e1OKzpg06+v8bpGVMgwxAKBQLRJLQ8Qc6cOy0jELEG
jwzHk9U5US6cLcZ7EyhN8l1Dj2Qi3DYZqAAIHdJN36qHy30Hk1ieY5q1KRDwmwQR
NOO8LeEreVX0vcoqsk+lVf5825VpyqSevO8SZ4M68m8MX/qp4w46vQ9vEDwt7c5g
olMNpExS4qyyaZxnUX4H4DSykBTc6GVB14WwytrTmIfsYndiV3P6dvIJdkLKhZ3T
js3Q4MbVJb9ymaiutoWI2izWApSgkQE+Vuf0jOPs4GXSTMlkbo5tjTE6wkWe+gqW
2i7CkSJ0ybS4PNWAUHYzxMZej11qwEvRDeQP7kuYdYcP/KrkFGzAo/Pof62MWMZD
ZdQdqdUCiUgFjJbhdYiZXJDa53SD/b9l6Cizx2nH517myOHni2Ex/T3HXvH0F9Ar
RuwRGNeEYxpBH6s2IjTyT1zLoF4KXRlFhZBfscyEiE0+WIWFSBogbh8vMPFDA2If
n0rcIuTa6zlMIhH4wKA7rN0oGHM/8gRglYNBKU9pkheTFt6AW/7uZHY4BDk4LFKW
n177qtsMcEY/oOBpgE4VTexbV/Q2XKcAgzey+m543PvhkO8HL7G88eerC/mJy3Lj
9FI7EW+8gNZIuF6VarRmIg1LbEz6GaEPOceRyk2c5um8C6s5Dfc4L2LaqiE6X2WI
SGGHZVftKasnSCvpP0Mridmw8EhmEYe3MkFWIHipi9SRYjVqJcB1U2WQC49Sbitd
fhRr70gkEJujUtmMsSgIh7tSElhR06i5gFzdbfDRDgt9/oeJ2YRPz+I0QlbMIdXZ
bJmA9YNu5C0r6fXE1YvAj+gyVRduiM4Pv4tgcuZ7VhUzABQpI7JTH2j0CcXUF8qd
KMMBuwfwl67wOton0dKn4qNfmlS5iG7XixjIIGCX2rEn7MfrtU5NRfF0jGqRUFcN
LA4Y5DZucHl4ff64re/R57VJbjr2fsU7G9/6PQqjRIuE0FIROCqG9tqL8ZqQcPHn
Ps2yvOK3WoqJjeFprWxv4J0RhX1LvjLBLTH95U1z1fzxMAaT+prVqq6oqslMCyVv
qjha4chkeeKfQSNZejMLkn9Yco0YdP0KDdkpDpJnWloQg7YlMpMp9+ClWeHVcUfC
glUc5UdXhP8ZKIYEeS7VcxZs4FiHN4/XAWP0mVdsqA5NPp2lkS49DK0s7CozIkq7
p5i1KrJ2LM4SOxK13fLr+irUHqPxxKft6X1/IOt/BpopYdWoEIBTD0ywNGfiDCAg
uBTMUcYct9aLQhgprvxObsWDKg6puScM2oGt/hoTUVPNwJN8FaWKgWbD6ZFYcMrm
3A1ptXmqEY5/lbdMIATkw1prX0Qi2oqaYCah3IIrnz/DJ37yZCmYUGbGQwxz4wFN
vT+8PRw1JgpcrA6zeZw51iK3uj8phW/fZeDDxlSwSrli+SsjWBOONYccY3dwRmZx
RKySjDd2Re5x/uci3tuztsSCUmcsYjLthKtk/TAmToiyD1tt0GWx1dtDxRczuM/r
bxEAOd92UWSkjFoBlmNLmfic/B69rcUueNtC3artyI7uuodwJlCiJlTYUbb47JYL
71nm0nM/ET6IrpjqmT0zFTgBnkV3jEtpeuuwiL/D3lnfmkayIbaIWN2S/G1YmEQ3
bFq7ZKN5mUS6WVebsj3xq2dntMhq6+Mke2KCyPO+gNb1aMpdyAeYzRujyUFlO6KC
Beh4jlLy1ZqET8hl56JasBO/fsnmeEBuKZtZ400BsOiEGpHAV9lcEfXSB06l79Ua
IlXmpOqpRJPavEFI/pvWNUCDholPQ/t8lbM5RIc9qTw=
`protect END_PROTECTED
