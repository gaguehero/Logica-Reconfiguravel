`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnZvHTAijxf+/0+XZtpJTpbJvCFUZNjtqTIZireEa8GLt4nyP8x2XefAetXyC1n/
glwGrSPupKvDwY5ruafcJss+0+Rp+cFbjozam1MFFxsn/IRuh7uAsCDvFnprtJlE
7JD38I4IyM4UabNFDaFNhEEevS1aFvgzbErBWzYWhryN6ii1Ec6mugSrWtlrU647
1l2VupAel+Sj+pOag24xT1ftc1QnermkRILQ7iWuweIggf/noEjgKL6CI5bKVCJO
gJn2E6W/A2H73akhzd+OmCVOG/GXZMkka2nWMNQqUPxYRfYEZ/CZQNu6LFskzPUT
aN5Sm7EUKaPESyspSF/Bqxb0ynpGxOXCC7qPB6A1GD5k7LCzOGA4yqlDMaQYUPVK
tdwXCkjN4hXYYL7hV/SUAfLKSBiA8fT1iqHHxaMkOum+gdfkcOWuwFJOXkdbihEi
nAEgID+A71iZbjY1A32UlGSP75y4IpErnnZmxqsLCz4GJIwg9f9XCUjVzqBHPHZU
PW8Lu1KiVnN3zP+plXdiGihTh8dp0rOnpw2sX2q1RwheNlJXa1y9FSBXLSuDFn/U
vpKPHunqVsrnDEGKNihUjX5IUGI+lq4r6yzUG4Js9UuwGneOhkQ92kLPdXDVJQUi
vLu/X/NVkPSaZSXl9YQ95XKP2yvTmx7sjgG2K414FXyBAUrzpCCFxGmGijCzIdj6
F34pkaaK/b9IWokAdkWDXQ6/nt8F8le4JHAh+P65pjWsLgwzM/UfK77NYh1WsAwM
ELa3vwsU2yRflzQ9ZHfMymwMIyVepX22qjGBGbLcvmUUzYQyY1FOGqCIy1P4oKJG
J31XJizvadx6zbSS4bfwt6M1YvVmzHWunCUuE2idojzX2mIz33EwzyBzRvHI8qEy
Ijg9uVcG7jiUYFxWrF39Pak50oltSMFvRq0I6VZqbd9LV0hYd92HKm5DXFu8YxsJ
AqV43HIMPJmw9GWb+4HGda6IffU3xcGa5ebGLjKsyKRe0Nf3/rl6z4wSZJdfOSMz
uoY6tlVBQufoDl/piepxzsLg9bCq82tgIBfq38SqeQuNFfduN5GzA2TWFF4pTuSl
Kmj7Od/wvxmlMeX8YSUwKnVpOCFg3J2yvsEtYMW9gAf7qoV11yNJAjh/8zzaXCUA
wPIqpY61zZmNe8Tyje4Ks1mR4xrP40CzncZ5O9wCH1B9jwIeoLncKdkM2SALJh7F
xntyuU8B9E+7QKxpbadTvGX/QoPySL28ve2wIXgUo06uuHMBdJY7qEZwMjlqkipF
/hMKfBEnQ/smCpu8Z8ZX97yWdJZ2huiuKIVrm/nKBBYkuy1ynxhZQuqUw8KdJ3hE
/wpbb1xPN9x0Q17GIr+JMldXVP8ItdISIH0CX7q728JHErNIQK9wckXJ8Xh70auU
xBWCXkf/sTscbCKk4Fc/WK7osfBpCdyXjKXL2dpRA03TZrqgTsPpBKuwsmb8zHtF
qRvnfBPvupq71Witt2qEBSiJcgj/xvcgkn8/OsNIRS1PJuSwTjHEksZ4iILsp/iQ
PNYicTiSgO13iUdnK448FOeeUXrxETHcshq46WF4i85Cy+R59WTW4re8yUrviQj1
70fWUx16vGM65W8ushgIsHD+aqWpvpld98DUo4TmkG1ri3yCvtkEK4Ii4quree4L
CSn8MHj19O9dnLfOZ3bPTjIJrVqkC1CC8m3fVFaLjMukzeoan8XO8Gq1xCGbjWx+
/tnWruXDgJVGTwy4S/Z49gEblnrCosd69UypZ63whOBuJk0j3v/6uqiCRB5ztxmU
qlNob3gXCjhYiLvGr3akmX2C70VMAo2aAQW6SisAbuTQKWo29NfmDPFljmuKf1Il
Gch+RzrvqohIjjqMXi3AjmoPTY5WsMitIgWOhhOpR1sdCHXVKlxURNduEKcWaC/2
V4KXnCrzl8afvV/16OdxOycrw9lwCIervXj2AGmjEVxmlbJ741Kw8amtSFsewiRU
uygyYA38hX08wYV0L2ROSBD8UuVtbTprykgpW3yg/ndiipF9qh++6rBsvXfcbmMX
66WMKMKUn0zMaibSVcHCOt9K//ceFDrBE19aJTTwOqhPPnMTcI04SwPutVdMIcLk
+8Hyfu1LbFHZO8n1uSoRORdO1KwTMsoX1uTLJmYmsizeefjGBQE4wYDtR52lNPoP
dJxh30jgu/Eu56tO+VgwMaFBKCuahkkx29c0rt2lUo4ey09LKF2DG0I8QqNLdXEr
FfMrWQmfew+80e/UUdzlW+CmA9MfbOWn4Ob4JsEWeohAOeEK5V1W6NMrzdi50V5+
otULI/PReyAUvNrke4A8Xf9/79UFljA/ZL2dSJHQnZwOA30A5nCbk5lXT1ioSxFd
n3BvZVI/SvIvaQi0O42OJC2zv0DZLucvrmELbmHvSYcp0Pklql0esva6N9nLRfPK
hBI5MJaaFKgM9gX//5A0GOS/1uW2UxyI3lDaqZfm5E8tWwYrWbsyzlIcRrl19ehX
0nnH2ySqcd6EA6RvfywOUZhOup2XqMWDoZwizbQGxSwXcKM+0nFVeOkRyPkY0vhY
JUnv2wq3xLiV6J9xjWwB0Eb3G17n0n5HnT2xNk02+893UIuuacQqOunZiVIx0tB7
uYwqCRysl/x87ZMPcnRX8U8RMyJsPcQe+ktFxAUdjrJN6DSuV4YA6oHuT+QbLpdl
vD3woA0CGlURYj0DJHGGNMQZvA3sgVfW/D+8gRD9QnOiaeZ7XHhbYU3BtPmPdvrV
k8AAdwy2D2l4kVz3rEsAECQaLmO1qKSmucJhyKQ74OysjlIfD2D6EY8iaUl7JvgA
+UUaxxVRlHiAPKsecLbRpqcQvF0egyvgCbm3m/2XLWgvUKI1axtyqiaWk/IQRDjo
8ujwIhzE8HYeKzIYuAKdmLnsowADmct16hzSS6Kz406Z5IsznMMyeYWNT248Q5yy
Ww0diJ6FcCMMz3RC4OltL2soe8XQVVsqWOSnWaUtwvnNAY/+SkshEnnljKLpBWy+
fljGkKWdUwLFIhcPZeZjsYOfC5NigxUldgvn5G/IFV5OkmofwyjLANzOYRj/ruHl
Jclgt4zuYxiUKK8lbIpk53Ckg0IDF6haESFJ0arohVdnVV234/dAehFIpF7Lq7/n
b0JYimu4vDSrFNnZnP1ft8bu1RuyqpHrx68hhqPuaPjMDwWEnUMmYkBHSQwAc+hj
GL658Q3WjCKmiT8lL5trRAIEIFcMuHqzUtb52e6PtWy1LsEwzX28iX8f7U65WFi0
2yMYpxFUrC4ONMKfm1DoVUm8+23nRIRpzE2v23WRnuqOWVrqmq4d3EJbPRRrR3QH
W6RCKn7wYPLBqvtZ3+PcOFEscxkO5NiHJr1XChuNqRNDL15DYdcVJDyhf6pQfcdf
W72nCujCIEQd6dKoZrrMFf/fLvGy/wOxvHHHr2iynYg53jvuWZoIoJLE+HqbgPtu
IXD0seA3Mg3Li5oVbwEYEOvBNMEEtpJyMwVuKNxG9Xtuo9rlf40Bjvn5Gkhl27yc
XIKS4h/wwoQWXTgAu0dvjCow4NiSpJqWVKbpEOukCP8sOr9nFcy3wPFvyrBkQ/K0
o99bxcjvO2J9piiunFkct/lQItfs16ybTP47HPLsBJZ3mhtF4i+JzjkRKDIK8wck
9HxyOo9oVhFr4iH0fVQbPZMvOXKj8s3aPMPXlhZ7iBBj2wHfC5P8Sht/7TdajgPE
Vb1PtPB2IiB41YFRvLXexwPN415rt1CHVPF5ojP2y1VB7WfWdX+KGZt3z2WRQuDA
i93mxYc+Dxl0bb8+Klk/NL3BB0zxTD3idjALJCGlnyFBIoMN5MGobHALMvnRPDx7
87qpEcNyPAQQAtI1cld3m7hqrt25P4h/M604oRjOOVBPyitR2SgPRPqhbk3OiADA
vtv8SQizrH+7+Pr2BPn9eo2kvMId+Uaf0d8ICK8Qn959SaN8QeYzanZCWQno98W6
iRq5oZUNjlEP+2IyY2lHpF1eps7c6uhpfTYDGGKV+Oq3AwROCjWGZ4qj3jKo/UoB
QSXOVLciS3FLPosMPdXYFf6snqySnZFBv3umxj4la4Cu1bTvcxUPygx88EMd1FS6
oub2OcUXoR1zKMwFIkK05JRBW8fVKQUhkfcvtE5yfQEh4U9HSqbS05lAdLIDMQt8
H25J/OrM2MJb1mUrBvivvMSfm+7IZ4NUZmdrRELi76QE00E8tVqGRmG9WdO4NRaM
K5ymOFxpAcV2Vop369LQHESq30zZArRiKwVVWno7WZKeDlkNwm/F1M9VVdBNN2Po
ynr/dba/ftiksJkpct7/7AHPKokYGmJxn4f6ETgd04fzDGr/bxM2CWDn0iKJsozf
cys7+xRafFhFomj6T9Mi6CWCdhaaXHBrBFQKegwc7UP3D0lrXlwWD6LrKubivcQR
KY1NX9HX1/D9QyC2CmBDqIKj5lYYraCss7dktjjUgtWVXrwKKR1Ou4iWFujd95Rj
60WjD4NjY2p4L0otIrgX/X6QmBk+IoNrsvIroviH0UjV+T27v/inDklExkd14a0A
NEYnAgut3YaYyI8Xz/Ph7FKcvYNM5+JCXoBipmHO1f823MmRZWei0M8yp0RTWuvM
vzTCGmvX/U2YVTp4ODjFF6usew93bL2b6bM7BffTmwMbVcPUOgyW8EkKW3wSBnkv
vuOSy/h3UIowA+XHfvEC923ktxcx7M5BETtES2pXmWQuLhQf0Mblh9Nk8tSaDnvV
Wxsnki8OFHMmYnlTktFaXcT36/3kPCat5OuZbouxzsVEHYGfoxzU1Rxvj2RBbu6O
D7QStzh2+mvn2FlbRDYjZ1x0rioaZDPVqEk9X+dziwa946zq4WLu0+Oy0vcAvTiN
3j1zMzNQO8CvIxXf25ijO00L3UBjUNFQtuPYUVWHW10adH7OpXNTPYiCOfB6C5Fn
4TfUAXgad3lJce+hyzPb0EtYV6be5BlOB06nFBiYm7liMhMqRO0Pa4l7zXXvZb7G
YwVjZI+9N+MSslTRf7p0meE3IAZkAoBBp+J1AWxtjK4H2e/Grced5R621KzCR4mf
vKxkc8W0IvP3nUljuVKOgIxSgyMx/VwepmoluCFEHPEl+QhmLLWI+49ECMnB/ISQ
5hr7zwUA7LMOiDCHoI8qonGYo2AfYoxp4zRrF5foFjmIM4gBDE+pw6Amw/YnPOVS
bhXpo9HyCxSgr4+OhIL9s/wsAYQZxNhq0s/1rfLfwrmPzANbDtWmiADLXhbqJ7DI
ZZ9gUQ6Uzrjyh0gB4qht2BTZxdIDRp2lUfu5AASXi27eytsXBg6I7Re8WVs8dDb2
9qL383NIKGQbJEx8crMVWRXMQKLADF3RoR1Qd1UTVxNtklovr8InBOBWs96MZa2L
kpvrpK7synMqHH+GTrnmPVzjE5C2u7F22k9BCVyufsfRzV+p7tEdZkBj5y2TvwOv
7dK+tupYKP5D94UvxpkUdE2/u5bZM7tsJvjzhaGD82VViBWSVx+eSktQT3opkyJp
3CtQk7mIPS1OP+VvxDVZpK51MpiHGkBKHIrzHTVc+e3916SBYmtrrpDH73vdwjzS
hJJlKdDTQCZFAcvYZD0SYbbV8B7mmhORAnZHfpP/WtwAYcZuMuZ00NcHjNQijvTn
kLpldeuPRt3gYYBcC6HckpTBqxqQ2VgHGHhD/vpKs/umicmhvaxW7lwLIIYsNv8/
YY375IjTPl2OXO0N5t1fnHHZUZF9kmpJ9rhy99I4uauv1sftH7TnKgFru73aLar0
v0XafjBzON5/RcD3mjhOHGGa5u60jM9IchTFrIAsCIlenhqpcbJw1/e6JQsN+9qr
g+KCXud1rMg11goNLiLDBwxJMQOcQtw7xEsIgU0hR9lOEX0Gj5tFOjCemYl5oyTf
YFxQzGpI66pZeGjm+TQs+zEArTJSBVifwiRSzBjCGF8y5koe/j8lrXWTVsCYkTQS
MzsLGapQsyQXObFV9rPqiYoCDgpPQTyBfzvMeaw87qLvIQVr5hK5p3012/rhZ4Q9
alaCvX/olqAQxGp6ysgmN0Z1BtgWsfxeAnvjogtYRakKAXNapu66jfJI0N8BcdwL
39vuT9pjjlWS9elqmMfiHO+Erd6gHR9dj5KbSOacXDCpMb5e+1ufrIvksnWowFrY
CBks+5wUGsOwJltuRzXNN26N4VY8DaG1YUbqSO3JGhzpqsOO6TQEQ647kR8ifaDz
8oqvYo2cNmZUOMoen+mgeymXf08nYUrpP/snf6VljtzsnEcDt9ljpcYEVlyNFoO0
QLIE7vs8fxDkcZ1/38nsIJAlqpxyaPLwPIlFU+JCrBgguAs1End0ltcxsKnvbqg2
ORIWGV1V4KsZ0DHTxz4Mo1oRjHVQbeiNuhdekrhjurbVUWWIt+JxRCV7bdbIn/pn
IselBMKBxU096nQo0AhYnYP6QQTUBzJKGy+GrDgKlTbSWiIBmDEfO2hY2N8w8qWX
Mu/LNUXGeQW/39iTRUq+5wJE6fYR7c2fwP/pLoSNSY3JQ39g+o9rjcO4pjdVUDx9
pcg1Qa8GoYZCS9hqIcbLAYKYWgnzj/2i26OOgQkxh/slgAoeraAmECQSWv5ZMl5R
3jBLxSArc+CHnjEdz7yotCEPXO+3oeYnA+3q+h6OSTPDXDSPJ/2Xj0w1tP+hFK5H
HbC7KV6u9bpVJC+F57KiXwkkrjR8XYGM/Tiv7js3IeMBFPo6OiJcgbfX8peY1gpK
y/v297eHla3Cghe14FhQA1vyZXmwiAVgkqJ+EeOZMWFYqloZawSYjWD9mc4mcNbn
skXyhzT/6W6W2YEGU6J5TYFwHC4IbREAKpFOF3N7Z79F/0Iqo+azZxT/gd6H7dQN
MTgyHWPHk+Hu25qewNVNS8YokuEV00UN1xuvZVQ+jHeLNF4HCoRuauW5Od19pZMY
9D7QIcgB1cEbfgXA2IHUr/U77NXaemtcRwLg7QwfYOkynnKSwIRbx6ZbBV/38Slh
G1arcZ/nvc9wLKaJNCxtHizabXf7dC+uvpdWRgrc9i9U+ZjO4bWAYeL+so2SScZj
nWo0Oj54Niqqz+aavMBH8CiNUC8VXjmTzDM3MpuShCX1UQ1/TxadTOVdMK57nQAu
XpT1giA/75pYg5xfv6tQtwD6TR7h2R5xczttyRbAoanOAQKBZWgCuNpnA4FwUhBg
f8+2bULqGYISqwFuQWZ3JWm7/9XgZbFijrE7RihMhUbz1PAGsdljThTXvA/Cn2qB
rpN70v8wrWncP1BwcbvnvQo+w9WsH4cd3VI3ZDk4Iq3nkOtYB98b19+R5SyqQFBz
C0bKZUH3JUVzijI3VUejjvO497aQ5N/kBF14M3/tN8RDZeJVb/e4YWIPn0eNiDKt
XZYKgIkS6pCNFwht+cZl9papHwLSjpxaLgsN7ngbcHLJyzyOZO9QEAIJstJ/tN02
8Aym/NMi9zoyalR4302C+rr3YSKtikIQ4XHOBFm027EV9HrT6no1+MPqPaflwvax
tw8gbShEikTBBwJm/gmftBmsO7rdhzLCKkNlSbGpC3wTJiiukohZ5hA7maLEzole
q3qcLNICMMoGYBkAjxZLNY4BQG8s5ekhAaWy7TGz7T/e5T22co50gzGa57FqZFSa
4x+gTdpoXOlnJnw1LJH6n4wZ/S2dBABqIk4MhkA0sZvmN0FjEDhkmI95Xmb6fBSK
4lffkXlfQKtKug3CORNY7A2hTdAXzCUOx/i+z7M/731a1mcJgXDDNfRW6a+IgG0O
6Mibl1jvqIc8YSs8bA5neBUWiU5pDMDGCGeIPKqBvLhLMqwEDn9PXzXKFoE1Ffq2
w2OruHuAGqie3iMNT+CFf5jCS3eWSvqDvHorUfQ/O41KpqCvSVtlMmCL+gZyBSpZ
Xg0UAXyFcHiW3Xb+xtj3tSNL7b4j+k2mZJObJX2LOFNZ3/TX6wkw1PswI9SYJ2r0
IyCOrpT99pNwHMcTxvGlLUBsDm7VeBfPNhKuGlubGXC6RaphAfbm6o8xmwSqlCSH
9/qmuqY6kyLZoFKrG92eKvleBPB7Qwhze0D1IzMHd6aqtzlPLrYzFepfPhAzoeOq
bJqrXl1XjxvNYbUM8SWswJbwacYAo+/eI6J3dNapnUBRyecXtIidTD71RK23ssph
O7wIV9tzQjDcPTfxGeyLM8d09NN3WpVfQjk0/RNN4G6+Tc9ITSoikrHdWQWjGUv6
222SUrKuFXYzQPaBy8QBR4W6Ufs9dJZ9szkD23zM/fq4r7SckZqbTjRalEkWDVIy
v+n7byWsWJIT/nFtD9ilGtBaNcvhDHLRn8lSriZTmtImfr0KKBxBwt0OwAp3JD/r
oZBocCwnS43rxPmkYVGYFcsBZOLak9twlGWuQLVrrPXXoSe29tTLmU6iZUHlWC+i
Hc30X+dcMU1ij4vptA2he7PuzulQtMar+h8w2/01unS+n29YD9Ll2RL1ilj90Ucy
n2qV1c5pevQU++GvV9P8hRRucQMPSwpunh/MLX37Ecrb3m8CBCqqxt8rtFSk49NY
G9DGDT8FvDueIBZtEucp/Zirj2o74SfQlYEQ4lh0luCmWYvAjRZGoOYtKZQvk51O
paqnDWCePGxMe+aKV3mwPpRnQeBgt4ZO1EmLujSKZ4yiuqbekocAPNXWjZFZ2NzC
9TgUkqNr4cF1oiht6yoxdz6Gp6/TaAx2HgD5N1+CzNWaDA6d1mORzgAN/LsYvvJL
pDJ0eqL7ftW9+wfqnAR59xQ99mzrd5W26hGJJH8THGQ/a0vEQgdi+PcNk6eoqIiB
4YKBtDyPCB2bJ8kdKlC8m8mPMZ61+3HjlOSSkSL6w1dsoKgf1KGxzuujeUmAd486
6YG4Fk+rafoTpNun6veunXQqcCdNGZjAmrofYWBCv/7mnb9oGCW0aFinmLlQtq+j
t7alEJRKyJaQOZNO/vdU81r4sx6aZdig/NAFcGbq6Kw=
`protect END_PROTECTED
