`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTAJ3PGdATWWB7boQwK6LRVYKUh5PvcXaC6t5/TsXg7Ej8lDSY83YIit5nTJ0r9D
+bbeONa3DDHHOtgEJ1r3US1oDcVsL9/S2s+jkua8o/f2DQkXUlVPbZF7BzGxG6Oo
vJ/xPpK7jWNi+aDaHq4LfBu88ttCvYn/ePMkJ36ABedfX/95nHbTaKxpgt9wyYHx
551jF9kdk6rHlUkMVMbhp/hJa80s+r2xLUMCBrvOLuMYAkc5EE9aVUzL9mkfeORO
ysA8RjGO8C1er0w7Nn4IdriuNCNWd6UU77BBRyC/AzFLgbXkEfcf48IWWGRyzFTK
8l1+ZfRGJqIAjn5ra3YhViz81eR67KFbyX15rH+ew78DK0M6A7usW6gWjljKCrG3
0bQL6STzl0gZml0XIvh6LFwrcIXNV0AGWmiw1qTAqnN/2IpsE+AUXhU6L3oRccjj
8IrHotcyTrI7HUlwRGJaD1Rq2WktOu6dVDCkmeedztBJj4O0WLgLM4JxMIhXkUNO
BTWO63Ug2j2/LfsD1t4gpBsupuwXDnzwxTnXgTeyTD6gJCdxWkcIpms4es9bxIe7
9eQ0mlI5jRQH0cG/W6x4KRWCJ05/s42PaTYZ3cNhX2lO1zNTgsaJYgrGwd7BdUHZ
5TSqyUHzxgatboSNxZeU+GAzuFal4vdRbreC/yAlVz9xmHyJgYaopf5nWajogQLu
qQfdM66XUOKzJdhfda9muOo3blNm1Gw1LKW+VcASIz91e/tmsoyK6/Q+HMHEBryz
s0/mvbjF9+sfA3iHMBgYt61hI70/ujBeGBkHSGrNSn9Falb108zrMHjy/FHBSztv
LnNsUjhiYtYuG0LCE3cOBUu2reiwI1Y5PnKOPbmO0IQR99WNiSbfxt/eaYMqIPX2
vHjsD8wrYDuro9urD+XxyZzQR/EQYfrhnMmFXEhj9W4frplxZZTccwHCC9KoSAAl
qM9Y1RvvWbJHaXUoG7lLs/VarJSzHHnFqKxy+9t+UzoqwcSXwcVQqEgr7yK20Q7i
Cy36BFe+tUUCfs7f2MOql8LeyOYjy/eVIaq4Gfm+YEs36aaZa8lXquBJymoUN7NT
XYeiVKE8bn2y2X9GxOifzw5iHtwQ4j6zh8M14kf1w75F+z8Uj5uYhXvgMeek2zXy
hdnQ/vK4bKerS722YSO3Y56FkQySDQz2JCVkTOE1JXMEt5UO6YYNpeuiX53QNDj4
Zl3Ynh2SKPKzt/ZUQp/eFRlx831mn9B3njPrgkuntfIwRHoxx//yiNzOFV2QKhzY
yPgRqcrpB+EWN2KpuJwSmbTISX9aYZs3yPsq41Q7A6T7DyCB8zIkAcGCTCwnlZ3K
fezbMi3gAuFfzp7+pJfxso7EIz/h1gGyJyG+ITIRMgMYvV+y746+QXyFDymJhDa2
L9f7dGjLrrEhZAvGGx/dv7zvcw12/a+m6ki1xDBVcuMxnOBvGEqh7w+CWvppjHjx
yGE4pCEunK5FGs9kFBo7mvoB3J1gIzJISRL9lS+3B07oDWSkUN/wLwM5npR5+ix7
kui7BJZtlnU5g940QVJtYf/6kMA8vWqO2/YTbQTgn0iytUfAH6Ll9NHTyalOI8zc
VpDmomguEzOR96R8WdlnEvMPY1qafunZC8m1GWmQLHTlP0yijUkXduQz1Q5Stq3s
1mXjTDfeAZ4zD4RKlps78xzQ6Qs/kE9ZjumqfHrnFAf8WAXrXe+JBXqEthNDm2NH
7iJTr4t++VJujW/hLISE6JcvkVXp/6gYmFrCB65QQkDRWnV5k/Wr3MLaZRhEOkl1
1UTOQdI8Pb+fcVR9yAgTNPtK4clEwd2H+tdWSO3KLV21evnWIygXvYo0donkniJH
pntNR1AIx+neqpOAdQ8HXRhDNEUuy1p04DQ/kBylqQxPsiuTA3i5drmJ+JRvtbJU
fJoqusp/9qOnH/G7oGSGNvougYZxR6En3anvpbOGhPKViQDPrT2Fv/P/vIlfqzwr
ZMA7l9LuZ/p7vps1hKV6QbYojvxzd/kFJ6uE+eAs3w47+yEIN7VuQAyItojS5JY1
WKIUSg8R4uCqjUtCsPzhfVQ9WupJeQtaKnKzNLgBQ3aQ0l1nCz8t1Sc/7/SaVTwG
IgeJ5dT6TTpAjk+vfK8U+gb66JVYGq3xzx0VCfW4SzpYArndBpcKpBb8Npm75ro1
xRKj7OcfZsLZZjTW3mwGtQWLOUxQXomgrsUK2rwWB8cYPfX1p0iRDkBfW0nXrj9U
qPVa2NBWNWKv2KqNgs0Jrw==
`protect END_PROTECTED
