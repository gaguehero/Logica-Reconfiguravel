`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7fOu3D9cEO9FbQVsxiGLBSdkZyj6jPG2Gj7OVdwPkfR+U8ojQaMDiRQX2WkIa2U
HE+rUA9C6lY9+C94xE9ncJQNIqxHNoA3UPmu29LeKfd/bktqKuECBqVFdEue1W0/
OKv5F1vd3ZDliR5un/EDIenS1wVYYYilDfMksFrYWPyj55wu112HPHKVaoe1f+ln
/k+jjFibwF+j5wMVVWlaLSbzE2hKT5u2YIgSYl8LtmwLSlFsAsQXAGaYBaFWsJ+w
NIiGDNe4EGMOzQygPIPCLdY6IQ2eT7O1ozHESnYeHU8h4mvPrRMXyp004bYA353R
ySHan6OIWcoZx/5Bu0UHO0h01VjNhqHtDT+h7nvxTJlAJurXFlQ3qVJU9uWOA0Li
uoMhwXylQJowtUpWlPzEwUF8VDPBx7HgKgAC1XkOEZQPDazWh9eUv05A+E6IUho2
v7hqmMimIFVmeomIsiKOhwm3bkoRZA835L5MNANOkH50/BgVkX6niUiwhQ1ha8Rk
VYhoBBe93dTDOz2eec6J7ApNtXQr8NRg7N4XmnmSU8o/03FvJ6WuUWttzoT+nq7H
PKnMJOOyf97/ya3AhXfvs+Xag2w7yh5TuXlU4yQ4MT0P41WaI/GFEB1z1aKdQyWI
A79hYTbhz2vwMiniKHsgsPe6vzOISAki5DLb6dso57HvLI2IL4AHfgQrfBdckF9G
mNu765DICATeUp4S1AzyoxOW+Z7dG9R2zq+YQW368TYiDQc/y0sMgCS8+UTwSIWX
1HzvrPEgNLnuzLitqHarbi+DumcdxmNaABRnRdJ0Pud+1aogpboSvVXVy13PpfIn
i/cbAib1bGcYvVAkLt3myzZnDGfrv8ery/jYo3Suv8EWhctS/mRPiHxfvOXmbsaL
ZAQu1iTSDvlAPFUhs2PzIN5XCfWai6XKP/F7j2npoOPNN3F652e88IYSj8jR/pUC
+yjSbXV+d4ldZ/0WWnxDufmHLbGNySmfeik/kf/mEhxYAZO3b/7UbVv1oh+0luXW
9TbTzhSDaufVgaM8CY1hzqwpSUWMrg+uQhQ4XrySE2+OM0BX/3Nu6S0BzkZ0ETAa
x9YorliiVotI1hbxq5MkEuPrbqJwl/9StqP9Xeu9I3uw0+DzAxzVRp1mgCatlOjk
VDC63TWQiVx9MDYfnRboP1JkyzFW/ol3OU5FzlaNFgXaQSv9Hwb8rHXQghbgVnnp
388JoSeyr5QulvDm01v+WlcqROqJ4MfcR3OKAjtnBZ29Yc4fRAZVlWSH7ulNvq74
R6l8rwPKE+wwXr4WUBi6cz8m1/xVrqMrj3AbFmkUq4O599xsl1ZTlOZI/wO/vuwi
RvEqmog7FWZRSuY2myOvJmeXRSu30cdNr5ksP3BDrQVk+P8+mD5pPNiX4kNXwb+q
7CJQAhFtnOB8XLpfv7aieiOIGlMkDE0t3qW3XwywxWcYCtY15XTU5IHP/yttDpHj
3lCCAlap53XUpCM/MJNunMll/7DqvH09clL9apsRWOn7/YPd32BQHCf77pNInO0i
GxL2xuoEEpkjQSLNx7StOSVCMVZQJQuCINdBzgo7Rr+9a34Qs42AcCaCLreiBev2
zPxFtdnj0ZWVn+EUqfhd4F/Fd5FU+bk5VO+0RH45N8c3obp14cc7/zXTAPhWuK/b
glXrvdmjfGNsgU65SA2exjKbF4LJxQebAP+vc5Cnc83qDbAr/KgIXKz3uhpaNvmL
slDzw/A+kW6WmkKvsOteFaAhwU34XmtU+p5RseCiDPj8NISxDlI1OflsDG5qFOBK
NXnvCtRTTIs6vtykQ2X0oK/+RR5GYsTX/CKhPqefoNa9ht1fmHktnPFDVg2JR3Zc
BNLZZWkhXXGwczLZ4OfpHMfm21ODEJnV2Kc0tdm4bsXgYeXzYZm05QtiwnKwV9y2
5EIDIA+Tcnieo1vO1cMAEgV5lMu+uQKLGP+WSlTiE0bCrv2mgIrvRQJkCxGbqQ7E
4QleaIGWISiyLb9yVG7+3P55/irTBtMsHyuZpgxGsmtHJjC0ShLpxDnHqyjw540Q
YrMum4MSmKHflDuvjawyA9oMEYV3hKadFMACxE3S3c5tSRxgJ04onYFYimbyYkov
YTZseo9Wbp3VU5HzB4cPTruumKEJfNUYnq/xaMBFv4GhUC43WHUFw7kQQZ2cT5si
iBQC10hk3Ym0qBMSyv06LbcqBk+QC+z2IOfIWTYh96winxlF/imfWd5pj08lzypQ
j/4wGGYy+Ip6bjQA9o/+JA==
`protect END_PROTECTED
