`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZOBbV+6rju8QwK9fFw9/NBhv5ZFzy35y0oquG6aEDomTz9rXki9b9CtK7V+TqFgz
h4PfjWVVlPPBoFvmPKncjmasaV5LFXUPBt4E5TF8FacrIkOBvyrF3Y1oqNt2WPET
4oYen1XU5LZWgOLMVTZaDYile9ZSjuRwuwhzMpRnH2CXCjoGAxFAqhX/KlapWZEh
nTM96ETnHxCupswO32nnuWa6b7av7UeL0YYuJNja4APXSa7LiRzyO7qelsJJZR5y
wRblehU36Axno4OsIAiQpEblCqHVj+kKkPlR+8XhCgMUv6DHb1EHeKp1Y8oUfeOu
aQs8NpQAB+0YtvWr8t47Y7B8s1aut9+3mD2zHx0nMRzurVrjgsGZFQ49hLwDrIe/
3CAa0qv5dcl6cxNZgc8Kpw+kMEGExfoXSFPhetq7anB70iV2J10GvHj9XUtdRqck
sFpbBv1gS+71EVscZlGNAbAciQ2KumInFRjnZiFukBtiBpInk9nqljequ2rYhz52
p2DAvvsaDgjeqi714g3SA2IbdxEdV5MUxYal48wA39aKUyXzZeKg+gQZaKf+jnic
kRpbGrxnYiK2XtsHIhS+Llt2p7LK2tu3IAJ4kJ/+O996Nn60mU21ODIfXkHOoizZ
ewTHW6Lg1FH481Fb8V0sfcVPxyUTRQGFlWYMCJ1t92QkTbCzbCreIxV/f6LW9ADT
OvqaTbj9ilh7w8PdBaiM1rcx9hJJxfnC8h9PiJKGK6cbT1hz9pcYohENdCrpcf+Q
8+nNsgo4rbunzHykBjzX/csNLVpKLcxjWQSB4jOuh09mp4docimp9KGPp8If3z3U
IMB2G+qA+4no4G6Bri0KI5kGcsc2PQqezt2lXVhBiExSdrr0KEddSFKU/q8LSc8O
XaKk08CYTXr0GgxzvKkDwssdyQrrFpLOBDj5vJw4Kk0TbrWotSorBij6UJnRl9la
jc2PHmn6+5b8yIGE1VXuUmDsji3DaeoXJ+mT8kYCP8XXjWwb19TfgN9IDugB8P2t
STjdtQbkrfOlddQMxd63pRddl6bZ9+COxWBTj3PGgeaL0NDUMRbte5UNlsZR31oq
6rV8QBbML9KxNX0IqNDn9gtUkyHdg5KVLnYBGUYl8wxDEJVObOYyRNdvN+osG5WF
GkPWYxrj483BdCObISawJ32GYtg1RydFFF2hKAwm9eamnd9zTjINwbT6n2cYmHDZ
rZxSwDb27qi5pN85bUHsOHY1b9fv06KXiuIybLeSloRKm5zLoLdl3MKpuyb+7cSW
clNHUTbgZ3i0JXYOkwEgoi/MpaEtyQtPseCiy6ZQT2Gg92hFPY534UiJcm1U6LrF
8wa1Mm6X9BZBrfkU6QXvtOdyUPyAtTgED9+71Y3SJhdD5CdU2L53ti7Gv6h99poa
hSnolKXWirx3XmQimZadbV+pLK7IEqyGuM9o1yRPKbPColcFgkks0wadJJwjMPDe
0SicGA2D22hiYjp9d5dBtXSkZq8wQ+OY1D7bx9Sbu6jB+htimCKil07WaPL0dadw
M7WgyFxAXRSK3B6Q/30QUiSf6cSe69J4YL3ubOcrwb87++hKJxGKZTTqSyzlWHj5
+JmqTVumwgVXiN5HdMdWvXbxv/VjL5bNUj0rIp/Xc1hse7egtzKO63ywRgP34ft0
Objkt+qQjdysdZW+J7fJveYm0TYYWD/dnR781AnRNL0/8qKLQaGe854tDnxWIPaW
amG7TUq/FU6g7fboXmHNoQgLu+Kcho/u4U6Z/DIw6KE62z1HbVEuT79WRDwj26nl
TcUIJb5TYj2p7HFZTT1dtfjt0S7Tfg61391Lh4ex2ttz7/Iqq79es2ozPf9OVMNL
vongcffOoZfUISExvduPbWor0W553t3kpB66QMcHM0w1h1mgVHuCYKbrWVPThiuu
86hqjYiqj+JLXXKR08vm7GwYte8Izc+vqc3KWDW1ZDNtPwbPYz/1iN6UzWR3tH5N
ewvCoWBd/ZMghjkRVpmpeyvJQaIg4J/hsPJIUW0aE9siKXHyOmTGsONsWHuQGv3W
ZpbDwwJLaIy1KIlPnua7Kfr/VXrdOOk7tiMILpY2Sevmgt84Tdb28dQnUfk8rc3v
3eqHf8GSm+gP4X7jCn/2036/w8WKCHJkjRqrQqPEyxdHwvV9cjx/jp7pUNnUwhTT
Av1j1oNVR8RzctiAriGe0sqkN2fdZiTuqNxSEoU4gL9lKp955B8UK/SkVV35oW3V
JC82Vf+nmxl6c3u4vGU5v445kzRGfCNCQvIHXj5rw+TotQxhFYWS30vSuOdx8k4e
i2sD47Dab25flh4QXIsK5s06SwDClfAv+KsE/tQOrFqlD10z9yBOUyXve3ruf/bH
tzaXepl8cAGtCElYD9pCev7YyiylpZ6C0ga6/PMTRP5Ez5RCXrZwQjgyq9U8xCRt
6ZCmki0uG0mhaeK4yxRoZVnyyNDNj15J8ookuk9TLGgZ25oa3GIPTNp4wqNB1fyg
lCMEmTjrtr+dP3Szz4xFdfm5Ddz3OW4wGakKlW+LBXa1ANogi8l7T+1ojS7cPcMX
7Cie6XGgoU0JjSm3Jr0sKy471yH0RVan8Vkx9qkrpa/GkioHRb7yR1QUG/UIAsYS
wf+ZjrzXIV/S81AwgOsmbQsuqXt/5yJL7jX4zuRRbwi08NQ8huKQO3BYWkes50Ys
LwgzJQLWOntN+nPiRlRF18r6sgguai6vG3dpIwSgombVATAIRc9IeS33+3GD0q0/
ap4N4eRagvYD9DpiZmEldZFxPM3NRE91XRbyojES5RxUjiY9bxG8vQAYZhn2HoDD
kl/4tk5v7yb95SNMuZlNczwNqIFhKOgJBwPJTYruaRGLGvr1iWAuUVuWEZ/F5e2z
3vuBjKxrOlLekWzzNhtrdFiiHriTMmwULj66DZKuVJXj98JS6SJkLUULesLMvziZ
hWpgbPgUhzfyJrnRwjSz7o64BqrUKLiKaMzM6p/nbBAbFexCai7z3kohzfEDkql5
xt6DCtUFeTSgAsF/gG9+ETxHgXdXDUkahGhQEe9wgqrIws1vJ6DdiufJCZIianMc
Nh5/6hCCxyCV5hTSxsMFNnO/y+02H0rdCaTL/ylUPk/jibnlwe5PpywUPmA/o2mD
tAEt9G25lzhpZ0clSMGsvVO7I3R5UGhU1KNtXmZZFNPPmwKmuw3bH4n/FIcz5K5c
yyFpuhQ2MJx7w4aoX0c4Dm48nqOi7ZUFbU+/57J3ISEQIRGbtkTzM3CNvGkzJnBS
v01brgsM2BhKrHaaHkFaH/AEo8b4cIQKq+L/PCr00qJjasi9JjsdoRsXRJUawMva
DscAAhM0BqFPuJtry6lvwHAE3ZJbBPNDlo7pK+LI9OPGDs7rj9faGqAOpuQVExEM
qHEWrZiyv4WMj+rikS6kDfofOVuNIaypD5pK1oDMmvQK2KHXjhTPDiUvLWGwfI6A
CIwCUuoG6VYTyfErqSXgdAaiRM+oJQQjs56VRilES92WL/aT5/CxBnOEfEhMb2/U
LJzkdiDD/7XF/SGvNBJEHJ626DC92c6Iok7FCPcwiuN3Ur3ZXU1TGJd1pltgByY1
89tHJnMrBuehGzmSFwEPQGb9C7UKOQfbvAmoiyQXq2J7GFyjjF2r0GwbfwyY40aK
6DKVLHhtUA3OX7kb0y0xktwE0JUf/I5mULAQ0bK6Ykfkus33T7zYkaaL9Hm/V9ju
+9Eck3tyHlqhRZhHDY5kxjz+9EqdhKIT8UlWA3ApDzFq2PdISw6aEHtnXSeoCEle
TNi+iNrDztlbQmOuA5kXOo9wBGSSIz40vrUa63oji+R6aupOngevweaPB50oSiSE
Ivh/yQHcOBjEofhLQcL6WahsnpQzSvg9esiGWYxvb2YL3aaUelGSbwOKTIvGIjAJ
dk+lssuGp5jk30lKTKRENzPDuo4zB7JbrgiLQVWFPDQtDAfWRPh2BtEUD6Iaw8Gq
J+OnASed7ey5JumaTV6RaAmI7jn00isq3q2cjhqPBAv8ny7eGxBWOa02BfuU1UBt
gkSKR8b43pyRWsC9ZoRhIwkYYtzEuunYX9Yhv7j6mU3gYiqMl3/n7KtyV8bzX9ix
KOi/2xQipIR889rIYFQOFWuebblQF1X7bcw79ZLfga0Spj04iwyVvQOqrJyQ8jtT
U4GfggoQ8Cezswp1uHH8VEHM3iUQ0rvoIkTme91f3buJoZg/lEp2c6V3fo26PyZ/
8HFQ30UXVf0DRaKGdkThRBs2MMBfElMWsRrdOjYZTPfwHivkGbMwygihVTpbLFDz
r9U00bMIPXvHb4iYXkExrazqUmzOeVNLWAtku3odJFPBm/CuyVKjbCxN+U/7Piq3
YO6TK4HiSrDHbJJiq6JMATTKpMpioXSgJLJ96DThmBIedbFgr9ptFUie/7idhOcI
CYXjNx3Psc5exc2yIVYL4qD7jQ0PIqjxG6JkSSEmsx9jncgTZSQ0D8b0gKzN5dvC
chdIIp7CRmMwL94HI+nzGT3up34732pbAHO0EcCTGyWN5nA97z+mB+BigkMGXjjG
GU5NDsonvXtVffiZv9CxsPWAHzEQo2nlxkhi+RZ4Pt0Ugag6ISH/2wiBaewPNAWt
x5BBpgGON0dykDQupgX7MaNvZLv5m0uCA/Pj7RPOEQT+egDOTqdJ14I4npQvbMg/
HhPD59k6kBkKc5xhN7okbIKC7YkPxsiYcZfxevG8yTsxGBz5ozQW8jAAT1HOcJCk
Vlt/ojXyCvxlDMJrNJdJ4DkJDE9a8RkMQJutQTnaPzCtPrxSf2PghVMkM0E4RX+m
EXtItNpuadL7Zur8WNqiy652chS6Nts4kZQB4kNxCw9yWCw1e+AnUSn/KRSrV9Jz
Ws9iogkChRzNB24PoS8Aay5oAPC7gQ9pg7isKJmmxjOYF0qHOOyZCyI8QJk4stiN
hgF/vDoest8uFi1qu09/6TBU+LP/E/bvs/M0FvkWu3qD2do9v88tf28a5BDS/Ltg
9mgI7C17cFmsl7BEJyDeCTLrVdK6N3ivMM+2oc7LAn6WXRL4EaV+RnNY3w76fPr5
PaOkjOAPXGjbb3TvdXEG4E0L4nFE1PBPYY7s0h2DUbhDaZ2lHxNL+okFj5jWTfFg
ZgTB9LbE7Sq4aG5QVKqdmqStjTuQx0qq7EnEW+tN0tcDCCOsZwA0wED81khQYsPR
QJfEuSU1P7ODdBPBck/LdNmoYdpU6SJ1kQE4ZwAsDtWkWLdXULaSqaRhB3dG7A3q
LYBxb8jTJ1EJNDJZtQ5HcfLg/xTU9z6nVrYkOPXOeLaCreWO4dHfj3JC8B9LGWlT
ddHIIVZumP9XgrNkErj6IzotFUVFaNs/A+nyPfLEYt9dLIM9loG1HCV1PfOo4vIV
MuPfnPhQ1Kw70rC6OFs9+2QY5F7prQJTVS1bcoCg7j6pnLsEo1a7+dnAqm0uV2m+
ahzWHYdwvTK1Si54sFjOZKbeGE3XodWURFmRUNyyXYOeGOxXJ8Yc9CFdnjkCRP7b
nyGvFVaJ4dIzkokDMmks4A==
`protect END_PROTECTED
