`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1Ib/jqNKgR6nWchReJhW8rEA6jKXs6KFuxQfHmuee46OkWTndD4VBKI0HJadSyC
Axwl//68pgYXucQrfNAY904PUfkVivgUvL5Pcphjv02RUYxDhSfu3dP7h1pkr20Q
fZznjSkgM4FyVSluHlk8rzbMp/ySmT7hXO+rlhpSXFKGdDDz+ciwgbgRBQXnk4O8
t+wwTI5DwjE38EFnBXcy0YeAZZiHk1MdKm8j2N5mU0oVOdN5eELw+OnbhQuljCUD
voMODqC+uo+cC/Sh7U+FyjkvK3xb4XAZDevSDbeqSj28VBE9yamN2sEBYOI2yRsL
XqYjpcLcC6tJIZfHt/e4zX9d2cLrksoO18wkFgjxMUUB/niE1VbGhFf8Sf5+A+lm
7rmKzDeveyhiqbylSK49xoa9efTQiWTS7FU92eBuQq+Tmfc3UmoIrZAUZcPzo8OC
SImXAK6BP0UofPz/8EHl5g6jlsOdZlnYFAoBH/HVOhwn1DG0nSQ261PQD0kXyjVi
UuWFCfgIXa5XXUBIQ2X9TySZU/9IWxZNqwXuwM56aMINWBybNTm4JN2caEXGb1Fe
31K9/kH7h9+KhPMIcAWuNICGAmnaFmj1pvvvLRGQKtBtuok+JEdU35a0u5MaEiZp
d6cAPV59W5S0icyyX/GA2mVKGXQn74qbT1+8bmkX8NRdLrroOtKaT4iGwHD7KmlC
ZCBcNfxmiViJEjrlTueMD+vJnFJz4l55+X6dZqca6ej/oLf6SjjxQKAcT1LKU263
tzkez2Ppi5/KtQNuvEXgpBjDisANEvWDFy6slPKlaxpJU7lAlhRUHkGrPFeslroc
pX8CqbQHvtBcH4k715MHvr/8EHvgLFRMmPHdMflrNWWtd1/F3Dr8mM9EP7nhUxY4
p6Mwln0z9wQmslnAfPfncGisut5VYDIzeGiGi8W8ze8OjpQsphW4SLaPdTgicRD2
+pvaNeJyxwZ/XaIqVSoW15SiSb8TKLCDf4KI17U9JGW39AtPIK0rqD495Ps4B25/
jzFxvC8AqvPXD9N0HWNvuoUAl/F5ewKiuC+Wk//LlLEkUQk0RyspqEVcrobZFapZ
GnD35axaEv3kMnRL0Fy5EuOvAezQSxQqSmhztdyylSK1hljyLQ8x9jChP7jjAKzv
rr2pic1P6PDhYr1IdQU5tW3R15bEhTi4YOWMJSb19WLyf8xrsjjVQgQBqT4kkcS4
LEc2ERfGoe1zILnQf74LFFFTsCRr5JftrV7FSbxNHQejYe0UlXm53j07xTr3CVmI
zt1JLnidhP68uxaRxiLWtUp0L3myaDh5bc/HJFlmZ+rYLZuTMVs+FCVmj3ZQ0B3M
DSEJ1OkS74VMWd7TaVcQ1AjVjmwNXwbK9pYsje+6PImXzFU6eDyIgyiPavj6UKCs
Yju6g6RFLbHgWuZarvnPLxzx64QDQ7QEqitL/jESCt01hpRHNioz2fd8mfFJYY5N
joGCe1GSd0jfCz0bBhjITeWZqGtOIv/20BCtre+/haI/JS08NBhcXjChr8kssDsS
EyQPbdyjvP4Y2pYuwkLBhg5Vj15sO4poOaL9F9WfqckD/BOlO7S2bymvhOewQuq1
mRnJqFNDBQ0cAex2V94VzCFPTpdkQ4b2GnfvpN9wsrWYGpasvqYx9bO4et8QIfe9
bpvvREduMpAJAwO98jzQMlZcSrb//Uc1srkECNqb/JxrlRXMr7sLYP5REHnDsZdH
rjp0fWD1p+cX4I7x/3H5uS/EmTh3U9iZkCld0JqG/tUnNjZA9ajbPwDuH12E8E9b
vSwsRdrV0PrarpdDm+b5LqK09gMUiM+e9NkSOt7AlbGBrJjd+4ZfoiOL7JiBnIgj
cIsbmd9esqAzTAqkeD5ql06SoxGa3ckvIkqf/7ph2Pe+qj8gvi7v1mXBmrL8LHKb
0yl6OklD2+ixNnguReovCGr3I5ZhzkhQMl3+pGOoee+frIhEkb0jCkgcqRWezZZr
+bVpMkRP5TpWUnPhLOqKfW/rDH0erLDbktJTvp8QiAFZmF/PjWefgggX0h0VMV06
X91rNOkpS62pnDnjOXfG6bRkgMqLFwvQrS3LbSiLMsu4nPE0yFCnBVnsFGf5k+lX
+jaQlB+dci7EUNVn4a9qpABvowDRVnTUkvGAdHR/XRlSfCVWS2AcDInTQtrpiJ6z
nWluX1wsH+h9VIAWD+Iv4CqrtPRP0kiOmS6qlS6hlc7XkuMhbjfGqbnI3E5Z+bmJ
rrJQRXEnhTegVzTHwfmqZPLjQ9+j6eCqlrFPU7UY8gF1PvSJNYRnjnevwoewHv+W
q6WIl20/Lot9PdKVWJ25IMNEvr2B24Wqnyw9l/MKmClUwVZ70YQFlIMDNoV4JOXF
K9MsVauzWQGBBQXgk+EhOSpF8LpPGNUwlkLxx62u39gekS81EWh9HReJz3idqAwT
aFt+/uyvLBKs/HRcxaeNfs5QTx6DlfY5sGeFExN5P2LW9DQZ1t9S3UqiWsQ86zUv
Ua6g5yMr1Bsv6xitA9jOcouXGYbP8v7jRUehvH6S00026FFdDCJ5NfaILQ9Xodkp
z5DF+oRLaxZCzrjE0/ILJi769hHx7YG4N/SeNEOfgk1bFEezDcLdxgsUGXjh8rXh
de+HLHoN5NEi2EeTIMSsZBlwOMdz1kne/LeEYHQbvgvVfTWIvAC5h6ndxj7yov1h
vLpvpzvh4t9h3ZIl83VW/AW+DFRIwS5eOxHCBvDw+0O2vqrZj3G3JmVEdAyUdfmF
QO9D2MVFwmvv57To/q/HkcFdgIrBJuKImWdWQ9zWLcbmJfWC9xDvMQJuhNCbF37D
nqIJAy7Uat0KnKipr/oaBLv/+n3p/FKywGScpkl8afycskba4phRGMF8PRtvl/KJ
a5TWAsAFYNd239+DZqtJQj5il5IIsCFAAOQC7SFZukPpruiKxaMKIbCy8vejVFKl
j4m1K3jQeArc9j8lVrHSZmXuf32WDNEcDqotWsRb9bZ4WpOExctLjbdwxm2BZfTC
ETJX5sPTwjkFEaM02qXjT5VQFSibahdHg3ThNFAsarf+KQMt/sTgC7ZnrpefkdKH
OL0wiJwpUDw6UXxqfUfSHlUbtsodalwF7L9APEfXMElWJoHmCMOtRn1ubie/fVli
uyCV1LqRYwEpz6ypLRsLkH7Qwo5xBZuxPMG5gej9jXJAhSq+0x7tyvvaQmt5h927
J1Y2YwAsf8u5MWvd0BgLPl7/BxaSWWWacDEIbWEw6+6qXzomZCaC4zCkp6tcnRKW
Q89uEYESYWcIc0x4566O69j9qdG1cCriubg2+KMVE0SDLh9vkVJcxAo7V0UonI1c
Onx2bZprjSutXhpI/ewCBOzaEfFdxlqj2Db+F3z2LafWx2Wyo8ujJDD5niKy50DK
Gqj8qfpMf51MiDMA/ZV+dqpApQb/0Fp7LSTlzb8c6YdKgn1Pk2SJppUrvLS6KdQm
IJqAD3bzBnTg7TImxFD3U9cpFYfqCMXNWuMlaRiEIvp/TKvF79OfG+xcDBMlDc6M
cK7mrY0ICaXK8Ve4SdhUhtWMGuhdvfOtgeX7J4wkADlDeVumU8pmeA/K7bRrqfst
g/X9UTjUqZk1HwxrAlaOx8pmwdBhtW4wfzIM2ExmsAryhyYyWyITpQvcwP/CBafW
f4b5nChyB4BUy17TyEJySmNpDUfxkc5Uyl6did/csgySQnDGtHAi1pzGGMQoZCp7
1MtgmJgrVAgWyjbgIWG19v5Co4YxUsWR5w7mz1yocKpgOfFkhAXeys1EPjVQ3Oyi
wA/UxKKZQfXp/3Y2pU7QXkKeczLgbdzoYF2hFHGWn+iu8XTgCAuHKbIGNrihLlJQ
bNSaHZGX1gaKy5DP+duFWEzlcJ5/ezvgMckthTQ7o6Y5kJ+8K51PPGh0pIH2ufOh
MoDXtwNc3rYlMI8okMuJPCchZC/imADz7QiaC5CtBfp7ZS88bRNHB5xmvzXBazLk
ttQIxI/f8ZNyiYWfWs4nk6HPuIUks78nTklbaONIxIBxxgfUOzTXmCUGk4/nYe2m
HNGAwrDWlicOOaMRnccJO2aA7EPkncyip/xNo0bSvTmqXjwN7rbMTwJkJoG72psH
5Xv+gu16NT2btHaciYI5yMROonkvRrVX8qSqHDW/2TTl9MQ8gudbFTcE6UyX8NvI
ZoDdUPv2mDayLSpOqLpN5+6uMwVsq6cD7vh10fG9e+p24w027hj+4Vx8A09XBQK9
YQPQuqlmwyTJYS+gzH+INo3NxHK7X7pLDRNGtnm4Ipw7fMyKrI1tlk8IcwKCGIpB
6tjszy5k1QxYCL1Dm/Tf/kCSP+X1QhhCH0HvGcVPzuMks95Z2yIuAg0L5K1Ffcdj
ryKJmArcS/Rn3N+EWnIHPI68PsLkNRqgoTD11FSU1NbU4vM6iexv65VNlhv96x9m
FLaibf52Yy0XbUr8ZOFzpdCVR9HhfylCZf/2fh8uvtf+jxVEJfKIMY3ueB/GGoMk
LfVj39JCf7ZOFMXzD8kMFO2IHlA+2D1Q9YBEb0VHgjebxOBxKyjVLiKoA8pUVJzQ
tz/IbSXUrghVGDtPIxrHem/H1jl1t7OkJa/+baRWGhydaNLu8SFUjrqdCKO7D+zf
ETB7BfkSLCgnbUrnaDdP185QcpDG71tLdsDuSCymip8kGd/W7QlarDcdBVAOMenc
oriUB7CKT+vGvMwKgMfcUJCkbKOiVQyX5QlbhZga+nJVARyNcH1N4rFZtht/F3Nu
6u157Ny0I2JeGXwSfupXBYW5TqtFGTI6u6Y7yrwh0iDxoMBydKbyXoO5M5we/hXA
vZzUnO4N/OQBedr/vPKkq95Q2despD8+138xVaWFEOf/KBLA9yIIhKcv3KTv0Clm
Q0nGRxe76qjxM5na12kLm8EPSNBguKFk1IimYhU7KlUA0+IFYUhMJnVkkUZoGOIk
PPyTzsTAdHmKrE96sG4o0cmeyL7oqDFuwdTM4MtTZHqvDZp+7et9LsADupC9vpNC
6LYgiQqaBQDU1xV8QaS/PB8ZtADaHd1NetOGcWHJJbuweOccbcXEve0Q8USpqPhV
nH8s8C6Cv8vzbBKRu9tdCDaCcPbdpL4faFBgaVuF+kwm3lgJ94fGV/VrqvF+UFsz
9meB9+g8gjZM31S1nOH28HzKtU75d1OYym9fQyy67RwAXKj4nLNf2DCocthA18hq
FasbeEeecGcF6l6x58guIq7yOQtum4DkrCoNouOC2dwhEDBjccCgMW9DvJ76Q0Kt
1R7o0+EVNNxVCBzbQQuSqeUwiEOX3k1ilo6runjuu300SeTZYMZYuKMOCApE+n65
ofat65HDdySlrM5wDB/YE1alRPMjF6qyYjcj+1JeY6MLNVHPLsEeZutLDoqNJEok
n7lj6wCYmPBkiQJ1NZ3zirkpYhu6Js+Fmvv0UvYCYjj/H+oBytYBVvPwYlFuQvTZ
bBf38JussB1t/1p00KbXHlbVGaubCsYmKWil5U/M8IOckqysWnfeVHy6IPyuxYFO
RChTWpWshVNS0xFkxjtQwogmxScsYc0tP+m0qEJNCX8JBUmflgnPwwNMcmxs/7M2
LbN4m9AAP0sgj8BAJ7hclQ5q3u0YPQH/lzxSlUxBanLi36VoMqwJK+v57HGBKNBl
4CZltNbItF1bISItIMAI3LoLBT/59R1m9mkPlADamOIJgtnFr0/YhIt5radQQJia
1Rdks53PMGMCc2CXMpGpIalAyYxAJrwu5PunHQnI44P48MepFWVp/uf3NnZphXiU
FJlFJoagPLj6pWjC8owjwvU1LtqCiiFLPONo0UgEFrWNEshv99lS4Wt5v0yqw9dl
E4NUt/A2Q7uWeybk8VLdgFJ6yQtduh4VY/t4k1G+ZACLa9UOp0ne7VHFL4/nsunn
H9AO7Hl4LaD6WRVbL2eNnuqAR1RAtbs9bDGN+7MEglmYnBbnd5/52r+1WtR5ZYAq
JuGGmV4LfaT6EIz0lfsHtc/WBReqFs67IxlWxpWY5MGj6ugC3onxd94hCva5ihEV
EmGoYyB5pGTm8cUA+PZPMmF/lD2quPrvi6T/r9EHqhQ=
`protect END_PROTECTED
