`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/iIjfZhENRJp1GaWrZnD7pKMbgvwnsJes+KEdfKCm6M+spV3BtG9PHVgtI5DZUz
ar2wFNzrXI6TJZG8jKXtcfdhlhGgWCw1/Ks/ZBWyiEbSWha/da8M14d6S/sDlwnS
u3F9KlD/hVee3fR9YMmY7OG16fGfYmz6MCAvJlwIug2LymutlZRIXp9MwmzOs62m
+ifP9pGqc557iUmcRLKiZucVUyScxVbX7U6MOhQdXUSCrszvcxjyzgbvBkWTTAhf
QThlVYUxey1FEZPlaTEpzrkFSKdEegvqokLFj6DkJfY0pl18MS35Q1MBiV3rsXwg
egrmQWDOcxzK84mcZnm0CCYDyxY80eziZxdIrH9KkFhm3J+wkVtH/dRQWzww8jwI
SQNMeuWVQs/vQJP7Ka8y/xTLO59HSyzvJzyS6IJw9VmxwwdKPpz2pH1cpZnz7bcS
leO8m26V4si1TTOnj+j61+hdgafsPZUS0o71NcTPvkwtuRVywmPbfJc7Ki+74KKC
hbsJJkpNjFVjvXd5EQhe0KVIu56slEfSexnMVENOzFgpHkYt27M+7aarJRTxfqs/
1Ju1x+4EmtbMatq7+oswbbz2uYrzCyw700OqJHqLreASmNeqf14cK4D7OdUADJre
IDK4Usqe2FZ/aKdPeFLukKKqDByHhoqnEZFXhQ3GJ8i5KrjDBSAdEd+uZ1iNsxQv
RQlbh+0JKblxc8aSpHO5o3lhivdnGrJjnGdkqwn80UJpDwp5VMKDXFyDV8x7BJic
d4rGZtMYDZkqIhOhYsB6iOkQT/TTo2Mm35MeKmj6Nc+ipZp7naiS3LLc6R8fyQjg
JvvPuCiS4/9waZbdzbRduVFh6SeUOA9c9yDJzUjrPpkyJZl8Q3UDq0gnuj9aIVwR
5i1N2DbFO9u9cZXdOKuzSiEhyvcD/6zeqWQlfNI3LUi5DmuqjXZ1vQN6OGVvp7/4
IUcEfthBjRGs8InoSOQlH4Lszvj95QF/zBYpGvJGJEIldSXZDvhIE2/pGVwSeWLj
Uunu3xSLOkaHrUHAvFOFwBENCta2s+IcZR42gdrhMzCjqXkmEZKad+JkN/lP0C3o
0ZY0Zo9rtMAO2YuzyFHFj8BBseB507C7DTXHg374kyAIpFUirQtO4Rtmj7WUTTa+
KXIdJmIcZWHY/S3qu1kJQSFK2dFzorDVaCOnsB+vg66OkVG6LNU1b7uJcn2Px/4r
YtHo28+2JYE5qtBjbbnBj1jwChL3cIgTpeS9ZyJ+4nLCcniHnL4SF4kat48N+48h
Njqzg3O3C2/ofTfaXViSv1nihtCoHbs85Orfv7fSNGXPVIVqNFTnFIQ3K+zYsnQ7
Nsoq+nyKpQ8pVIbGoshtw+DNmNvaNY6aN1StMfqz4RWafIAlzmRo8ErwSk/Pl8Xj
Ckewsk+gE1x9SCAsc2WYd2WF2TV6dgvaBxBZ54vkYeCEiDC3ILtmBxZz6Ka+krd1
P+zIA0JY7VjnqScATfqay+2PWERsFigx2WbmEEjd6UcRgwV4myyjh2qRuh7Q66X/
xlc2/rhDK/AKyIPQXye3x7vXYbQkgV0hYSo49rvGIpip947Q8datONlOtO8JvXt2
Qa4z29LHXuFaRzQyNZMiMedjDMU0DB2FHc8nZnohUcwxtzTBIqDm3EbO4EsjmpFo
16EnylN90c/xV31dKEQg42pkdgrpBGdGkHELfQdEqcEMbCzMf4reGvz0Y3lNJuEt
+N2HvlL3Eo9B9Pi9gJ2LPzLT36nISLKrYPchrn/DJtcamoZTti6RcWii5zy4Y7Ln
fbAqTsGtZxopH7m7MvVifIE3F6Nq8gRlHDH7FOKfrsCuFBZ/aljzFowYfhbkOxpl
4BcgeUfVwI31LWdIekyiyXWWrjN97635/zyOeANLUCBWlT88jPIpxhvoPNJRq5bb
3SDAHsXM7IkxGYjgsRCAaaRNWaoMkLsveT1hdlU0UaXhptE65e9pmgYRpOxAoi5H
SQNEXgHjGfK6WwJpqwRwfpJolz+S+0lR4n9J7MkYhVGPWHzWorVeFdYClP1ig7ba
Lxp5pEgnH9E81VGiza1Is7kARXMALtXSISo6mcl59bitD+9ciAc4DFa3D/ZiF/g/
6Z1flOG/cyPWRoN7F1yST70u96Y/SxJUcW+SRIM/ZCrG69Jar9Tow+V9lVeYcWaf
vzydWVzdibZm9BuGHCf1C1oTM0FP85H8CpJ5kme+qWg/ZBsDpEJ0xG4Pj01CGbzc
yQZN5NwgGKSkePpgjs5lo1MTvFxKknjOu+L+HGT5pF4nj4Bo9la9ZuiJe/MF57VP
mKqbn/9HSq/3091YOSFIMKuIgmZdvp0RV6AlQVkrFbZZmDE+mqAgM6xDh2gafvqS
f15/UxF8I3Y+l/MW+HSeMXlxCU+VbiGhjziqgv5E19OHrfBc+BahzXTQlTZdcJBe
o12A/45GGqyu9iD30V/6t3n7HmROmJrIpmRr7Zf60673cYUH8oitAM62eSX+JZo+
mOv7oyCH7H5Mh/Qw3aiw27VT/CPo/b5RZC1XUX8NeRVl79+PLHkBaYh43o/B8hlX
pfc0vfIqwQoW5P4QPA7ZWOH7S7U4ZAItiAa8qmrzqZnKTJVxzrPTKfxBxZTJQ9g6
I5zUqxMJa0VGsoZjv6ZpQyzMbchcGu8vUnq+ddAQeZmKynPH4/stWI09gRweoGco
yrIYJzwDvC/CIZ+1uhvEe6m0VlIRL17F8fSBN49iL8NZn+xjTWtZWoSA5727/gsn
DQ1u+rbFyFfBZjcq+Is8MpBRPWuNOtxKiUXHjTIQlWHwRT8ITD0Hq2NOzwr5bQkI
P+JWhWUwbF9Sfz4LWv34LTUgxUWe0SnAhvXzUeTLPtL4ZQQuEKh31Sc+ja82vYOQ
uBjxLuVpoY/iMmYfpntp5Td2Zhhm1+s6hxHgFQ/h3t7MtDb64bTyv5Jl5aSyw+TK
gA1btsjUTHtDKH/DlKAI+C67iomopC4MrMIKm109TEljaHC73ycyC7AbBvxz1IRN
uZKl3GF7dIKKfHhQOfCnbvQJAgGCACA/UuthJSb9H35X7k16RWikARB6Kt4YmeSc
KtReXuYaNrGPw/hRFAEvICN4L8CI0OJ0TxIYeK0Rd4bMwB8F8+H1Y0zXNln9lfG7
43KlP9vm4c24sOTmtJ+ML+9Zr+1Yen7xXB7ssVqTSCh3en3SO5V5fvID0v/kVPmt
3IIvJrcu8CkYFSogPItcCa6pV9nAazZS7lNZs79V098XfBp9oVSXnC2F0gA4/gY2
f4OYksgZAuPZFDfRxk+Gv6zjlMFvISlXN+3ROp9WjiUhSWeBRN1elBRXcNOrR1Gj
Ml8vDAnzdAynF21MOndsMoZEy3jMflb54GJdLjo8EP1EshIY8yTWSe+axMgrTBaC
N8OyESZQ8hVod56jKFrIkbUYq6DRNRx0uG+oR/JX+xoBH7qGevPThHyjtlvxsiTK
VSZvkwkWfI6yqb8CvAcbOUzoUvLKnaMMsZecMRRepie4cd5kgOMPZS/Hpy3QOjUS
jRcSkg+MTiitYZmx6grChlKMxBR4UrBy2ROLJATkld68N8EYfIgWvlnBxj4ZS5wi
wpH7g5OYtOr7GdKgtxCgcoYOaN8V3wxZGvswdtQFx467tX5m/L4uqOkGyv6iDgA/
3rWNzFa6M2E1DXnzvI/1L9IX1adxwJIUIFnZWUMVvVs6gUWLs+/0euSN2WI/U9gW
224bRix6wIxyF4C5h4U5Bp4d6rxTSWtds69wEZV8Vy7BrOalfYc2G+9PQTG8jc0x
aHyoW6sM4fgOf1OGcDZQC/JTfVryLjAtpFZ6WgRYvxC/1RkdEhdJwTeiI0VGL+if
UAxe4hFq4C8NVvRmb8z+sDoxzQ+XOUdxAXxD9BGuOkPc9CuyNYxXxJ05YJxixPfL
/OGbqmL/ErQf8oJF+64T+WxmrosXMHuLPEkRZJ+qDJqHoEup/4FJJaLDAyTjWY1g
7Z6UxBmcOHbl1ahc5jKbb4JIuGx60qEyqeKeLB5z4SyI6TOoUtKRoieipWZf1d5/
W4aVsIm+wRDG6TV8L1nQ8OkJZHCg6XRpHyf0AI4EDwXJMEm/kAMZnw+u0t4GICro
CAeZJGNsjuqa1gTetoZuGiDe5/GzxdCUwvCyUL+RTqNCcaPyUNGQ/tzc5ywpql3C
02vsA6w9s63c9d6SNzQnkbWN9kwZV9i22C83x1+WLgrx046KjqnOAZ4OQ9XyO5h0
2KLH7z45kYsp2nz7oIFOQ/kaNNP506jGUkug8KCwjV+Q7t3yymT2112/6krNbC6b
MnKgOyWJa07EKruwcFtiVxFZ2yh+IyQonXNSl3Wh0bnpFgQvBBzNihK4RzPThV8J
xVQ1rQrwV7FO69r3H5+iae8g8fV1/AKmGliXYcYTua8YPVDZD4ZWPxLMmz44K+m4
8YY1rriBHdMYXZrd7OHzw2ukSD+PIRwwu9a1rYoInOJd05H7NcUfzkPbaYshmUGF
zDfQfLx+AUb6UuxAUrf3lXWhTV7V7Qua/59AAXQgz7k1UJl9ufW5zOZ27W447PFe
8+988P1l09y9rmoMp75NfLZDgmoVvU3ooWS0sFkoI38+GSbdGcONz7iSilpW6tpY
VhwnsXU8eDaBgiu5PdSRaDoWPvQPZbQtHujm9UKWNAJ7b/1NQPugVXh+LimopRH8
MbBo2+syeDQmwkJyn8ZxclcV4NvSOiQmYYspqQoVUfKBcTfmSkUf1SfbJaTTKC51
9KpmORFmNU1J5VrGswJzdbZOwz3EKB9jzUv3rQWyHHKIzDb1zl7g3bfz6rex/2Me
rCJQd6KpRQu+MGV2WOwbEvle8Fxi4I9iQKwCVpdfSChf+/teQ9On2vvJI447IyE2
0HxhUrRfRjVNrHV/cN+fGivIo1LZ4HUwYBJqhxiA1Jiau0gimKk0h5yv7o3H7y0s
57K4/ZbCxUTTAhOdFltq9ATcJEeE/HFij4WbnZzKw3ePcdBjOZ0BbIYIZlzew0S8
JhSY5tqa+RQnMx6rvk+nDtgGhFPPVzp5Bq/bw5bkovDJKLVEms9kiuj2DgfwDEcO
PmY14prUjDbqBFqYtfRtq0kkBE20v4oJy4E/9B64dCbKx92eIg9Px3xNiRCuqiiP
YFDxPwEjcPKNLmu/yhVDWYekWMTX8VOoTddJ8q2HaIf31w7843LgC0SjHCuI7S9V
aB3eZw8nhzUpTYBaKvlhKvJRY08G0iZ0y3ZZgt3A+9bCvFFdgLZnz1+3E56zLx1P
+7A6fi77/z05HRZMKFpRMi9zvwxlf+RvOeudgyYPbv1M3cSiaafp4rzUaRWwvMC9
dxmiZtCRYJ637kRST0lGry2Cu6oqn3joechzkMYbUJw8PehtLV4FZb48Y+fNwAhH
t3uouwtQW7k0YbcuJ9rWzhXptU6f0aapqZc3E6zxVLhwOqa27XBvMagdRZm2O22/
HoazFmuMmmiO++FgowZ5icklSg0YGwLk38MP+4njmsFGxOIRYbJuhLVvOFi8LfDE
Ko8nmT9Lq7pfytVFgLbNAQBZyW+ZgVeYwSpWSsqpv4vdzSqZNQgpv8aIp1j/2xMU
ZI6Y03Su9PKZutCYZ7CzgL+NOh4291sgyACngHXYzztifu3zqc3R7ZvSNLqxFTZ6
6vAkThDN2rcW8vb3GeP0M0vsnKsRF9h7NxYG0WI13rJ4sLwaa3gO4TAvTGQgltK6
aVgVNNpYNgsOj2lNu4w/WjrMksEN1FdbT5IuMdyb9Uh7QcUl7V8naRapCot/PXKs
jHuMvSGZUlzZk23Gj8NKVXLB96X21Mlcy3/BANw+KkHVErg3+3gQkHTAetPnNbpn
tuPZ2VLYLoGdglVvxfcUoVgS0iTpZplhX4+r/nXOP2639wnmOM02zuzOORV8i8oW
b0X8q+msUWOKwLpV4BwRGbFAXaN4onYXTgXi4vHwPaWYgC5tDIdXZIjRWSz2viqH
xvHuNJjLJkTkGaa+wHw2XCJYWo6qk2v2o4VXAeav6e6prFpKd0dVq29mBRWH31M1
G0bC2/ZS185wAIIIJiMXFBk7hzYd7ETPRhYBqY/6xgr8X/jU5nZh3E90qpHZVoCU
grMjIN4Xmp5ZLRA86ck2ONu94t+3IuJmmj+hix1BJ8NuS6qM/SUoR88s0miHcQEe
FGmr79J5z/iNExMcH0zSjOAASXHMy7dLR4dimAfYVf5pI03d/lHpK0DQO5+xzz7M
XWAlv92B28tA4HkKXR7h+A7kV9qBI6vsibvNXvVv/8EykJTWLe3W2SVkprE8oh7v
yD3o2z7TnKRpSdCiRhrhQhxbaJFzVHJJN9m6ctv8tOwi0tYvNah+RyfpoKsvbMq6
C+p1+BTulYXyinF3D5Ln2oM7Tkr1RTIM2Wa7U1EzjUejVSSFYS/6YKZUw3auoWeM
qDAeJqTgWU1TScLNx3XPETsT3wniAspPKly5p2B6yyCiEnk9xH1D9wJCrZuDb8LS
XNtrJepnSLnvROqRpT6aY1Aowj5oLNG+kG87OuXDs7O33pljUxxpePWXzjI7BZ8R
Qu7qwElj1m4YRse2dSLjeLdfbC+O5UbVKaNGolfKBMW48XoBc0lUu93+t6WxSLag
cPXZ526+NUX28yZOT8cGUNf1GhieRdtCQM2mDvdnDRXIJbj1gtDvlZdgX6KhTWgQ
g/rVlHpZkjOaZ7zusBmhfpR64h4DGUyliBHH2H3Rioo=
`protect END_PROTECTED
