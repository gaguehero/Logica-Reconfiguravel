`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TiAFcoJdRnhgCpJKAMhRghC9zRpCaWg4TKn4OAaI5j2noBgB6U69v5VsRnOVci7o
jUBoZmKexnGEnNTlgzRiAs0/9oO/Si0Y1Y/3ZuCXYxrhBXBPVTiHjXhtjLH1Op7C
BCG8uifoNipisayCnIHewbd8GfftfTN3Nnm0Sh0hLHqwgPKUyYT58QiG6dPTs3nc
U/p/5LSIUilUg85cl84/o35OTM74wuuZk5gtDRrddeFA4JE78CeDHtKiXb5Eed7l
d2y4KlTVdSpMav5FTZmCo2ALot3e7N/4P8b8sSHZF5S2CQc+Go1JNuqA6lOK5XmZ
wOIW739DkU65P+6zLIIb0br6Ylkj3nx4/25PMCFOq1o1Hxd+013UIW6YqmRLISTy
pZDDXMNJiG+zfLscapDZN4OZb7LN4Lkw0AVH+yKBdm65AxXuvvQOX/WqHSgLlXWI
Ey/pvHZAprPArrY23CmJkqu3aLXlqPhh7N9q24OIB/SV9bnnPDLjAqu8VFxDI5OK
0YeENEUzdfe3Z6Keni4Dk0U6oGtwShW2kL37YVcBA/f07QciobaRrqyMofXUDuCS
fhPhKGZvJ3wowQUD3j2kXzTzOV2fmS1d7NGzMuq+LSoi0dk3Plk8y8dVW9Jb1Zvs
qVB4QJB9K9w+86esZesYj3WHpAgRBBS91HZdU8WqnuYqz26SKLse8liRC3Tp3d0y
WRmyjkDwiURJJ/8PO4cxHxADT6lbg1ZjrOK6Vu3ECBHrxCyB+sAof2lFQq5ocKAl
uyTOrgjIKcmoL/LRe25gaNV59TjO+wleC9ls2uP58WAIb5pzu+pMm3gbSkc6thmG
SEmnK5pasMiFv18janIkPgWecuOIUKzwnwdRuRQeCfd5RUqcfh1Cv3s/LVvr0dGz
6NsZeMilV9w8ka3FELiOYu9O9tpyQfS39NyNFftRo+M6T87IEHiDeT78ycpDEK3h
i1EMZ7OG3BNjwnxrPNMlNfp/2ozX0fFFO3d3ha7RZiL8jlBjmS9j3PHDdqHNybye
9efClVWo0K7shqSzSjOTich0da4Q8v/fPz0XVZWg75WdTsqyUVaJRnWJjnyx7ANj
zn6X+n1KsST3+YmV7fW56mpFa/ONUWYyviYnjoyQzn1rGlwgS/uY8NSPbtSWu5XW
6+5w1e/+nAyCNS9jDulB5/cJ6UYzzgBk4rH31mzA4bpl2lFWfoLX1QRGf3JMxS51
VOBqSOtpyKyuDnAbcBvOUDRned2R3CuCvJIjrW5dWoVxGbrQULwD0UmwzxmbRPQS
P8PjmT/rwyfwKqY0Ac8jemG04mu3G9v6gUbiAZkBj+y7bt0mJkeubZwQMB6V3zhG
QnwD/atQwMA7gnRTh4IkyZb2sSfgOPl3MxmcLM9u12j1miPSj9CaPZgPK+hOcGC3
JcA1ehPz9rBZpI5Q/RTB8i2eIDaPgBjGJdgZymLPjIHXVVir2scUMcrkayzdsGap
hcn0/q7Q+V/gi50WGyrDCEgbgVMKT5ytDFbFt0WdwaTkD4C6esXiHVho0Qz6zpfD
DizKPfrM7pfoP1D9AocX9kqAbWMi5ud2LsDeWH0zuamzU6JMraXHcehC3cdv9EzO
1GO9Q5E1NOjx09/ZM9Y6KaHvmQUrHpaOaCqHwhYuC0xZwClf2rN0sF1uuSu+jibr
QqVODZ2vGJZpbyjV8/1inIY6nqN27rsXdo//rVJGFzpI9jIC4f5KEfiT0WCMn4NX
rNz7064M66lf5u2oYNcxE82mvmCutmn/RWuEeicvUCdKFkTaKHVEHQyXT5XxBudY
E1Rgt+MGshS/hQ19fEGhQTU6vUnXyj3IgL92469bQzm3gtGL2p6mmJm89LuovVTh
/r1zujEaQnge+tDLIFdJ0H8dE9a7BhNW3/6Xkh8LHA10d4ZxmPXexUECmlLywtEN
kk+ozSAXlwvbXU9hTKQfdZWUwOumAh28y2rVhmBsCWVKXeEeWj9PWjj1JkQ0mwLa
JqbymSyXD6sWIIVNr/TUiCqEG1n1Zxypi0k+/K1FszWQFF+sOOBdqqvmG/i10xgt
`protect END_PROTECTED
