`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyaALg0wYep/FL4fw7Jby3QSs5CqcZ53YIuCX+8mQv+zF1jqZ+mmmfmbywb2XQ1X
eEybRrYJCJ5KgWuQ1q/BZy7wz4UXe5GuiFPi0wL6yjBhSzzQoNGeVFMwFHo09VqS
ODO/isx+aWTWiOcsrxFB8n3CtegOFV6RKAMry0dJUSvw1o4u1/D4/LGwVCvmq5C6
ik7jGn4NOR0zfCeAOmc5GXsAbxk8y3df/toASQsblUuQcJZuJqRt+wh7Wb9dYlM2
VE6NejdaEHCYwN1holoMBgyK2J9MMQhqpXRQwKKpgyhTM8GV/lx/6s5yWwd4AkE3
g4h+EHN7ChglCnAjez38MEa9LvHdRtWlE1fnBm8g3j2cxZ8dlhTGmLNQ6ydIaqk9
cqarCfJk71b7owJqSja0yemZopoXbUsv+A91s2P/1f0aB/y/2DRJXn1pxEPWp4xw
VuV2u+m2dJSnyxL0IBXVHV32T1oQ/gLMmrmJVEHs4PnY2Zg+pzYIHc17I/uiyJC2
726Z2zDGheNBNdiNV8iWINbZV4e3jbuiufdwuCyHfbok/KpYCDpcVgSnW5XPp1C2
/RSysmaK/fpKxNId3C6vOMgC5tInFoekSRudeSGixRdO0Kn9QG8yhjB/fX1KDG2T
cUHrBYe5TRSDb80+DFYy1IUz+drs5KRThODO/io154I21W7ZI04vz1YLSvbBILTA
j/fK0o5FYnbeC/cL6/DJ3Coaz5cSTLC9Yx4bjclt7X/6e6ZYnL/Vd0UKxI1X8TiC
RseCW+SKQk4UdPfhP0HgaEU8qE+sE5P1sJD72AP7s7Mte4hT+Hp2PMtsUWiv4u8b
JjQVrQJUfiqK3k1rP8nqFVmh3mb90J8We41KcRXiizzCHksCXqb5ZyP1ktODwrN9
nlhVvNZBXgPm5pRld2TlibcoD328bBaYJEWfeY/XhwPfLhTbTXzHkWLcFYoqAlVp
5sP0UWJPvXk3kla0iqSy5MFqIxOiqesTJFT1hvqyaJVKOlqUfQrxnWOyHdHa9UaY
vijjhmxb+xFFNxKAjfYj5A3GUrZs+WWyA+R+81stsZjBJFGe3dofoOvPuChIByMo
VdAjRH/SsBygU0XhBF8gi5zwElkD0NrMdrbyq6PMfJZH5xXnNYBkLaHuQUr4PHGz
eCChCHr8YFvm7e3iTPPtLI3HIOaP9FoW5TEQGuqYAwDMbCJ22/DRqPL6qtiXRtrB
3eOBfzty9XzLGrNr+M5IjqQi5/taJVQks8vjjorXhdWe0ZLX7Nc/3XemuGTTvTKe
aCUr3qk5Hl8goDMek/QuhXoGrEoDqjjVkSoWGaPdnpNeB6lvkaYQc4scSeoGJ0yV
nmuwRKh+7II/gldkMehvCKKTiqrzQNVQ6ULodnKYEbXGldTckd7ANg/TgVALOMT8
iN2JTLQvyAWzACe3zdjBrKIm9qUTPVN8G/I9M5FOhhsP2Eb2A6PgIxGwNBDROaFx
5iaCwBe1M5g84mS4UUuVJZ/XKtjLmot3/0jWR09Z6PGVTsdj8v589TmOF5UdvzS5
WM9yu3ohGypsyPfg1vraVzR0sXMaaC+OWSizfRWccpMNM3tKXn0kQgjCAfv3fcPm
x5G2bgunQzbEjZGLd8Bp4o9j4/bx2mWNupMOOJr53s+SYd3kCPlFqcrN01CyYeH8
xHr3x+CytEV9i6gXkTzPbuiIzmJdwwCUqJxchDDWdyLe7kwe7fwqd1v/eSGNiBwq
0vzBdKFvpWSr1F4esv2uipQiZf/3gqa4r/anp/Kld0En/IKeJq/ZQCpsUKqpq87N
8VmqPWPncb+UBpHIUBw7dtslXKFoMQc+UDgfxbVJEKG1HEDEKGHX1+dTn5YamU41
PaUe9eFxxEIIBUe64rKHsX6Ep+IzGwRnU+xFZQa/2dKR+cp2aVavqIHJoPr1LmZO
x300vdJYwqjyCmW/sVz5iP4aB++hn7UKps2XGPoMIfpeohtglh95/BOmf6ndwRgE
GjM2/cBE5mFFSWCQxvyGpd5pMg0zSz+tzO/Y09IKHVlF/QJDO4WrJY6TQSVkbFGO
gRjingvvaRyusL0uvVK1NUMVYD8cy35J6kPXgiWXmjulchO9sklFA0zpgFX6pK3O
fNgAjbzERnr0InsB59oN718adJXIlJ1UaQhypw/HDMNKmhtzYXtrm6Qyqpd0Fukh
uUlNs2cIZwLkdQ/tSmVUOv2Q2dpB4P8cyC7FiMo36D3vy//gb6zt1kUG54hL6TxQ
SYOB5kSsJ65TP31JRjN8oA==
`protect END_PROTECTED
