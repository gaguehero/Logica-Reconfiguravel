`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ly9RqiFJJYeD4Eii4T4Un2JomSgVCkP6fFo+N5SO9oA6uxC15zCjh+04lZssROx4
GfgVapYSf/0fIoNrKfT1s6zkxPNa60LMBN3FO7sW1xpTkrvYEgWDDcDLsK9m2Hq9
NJ8jVskf4mRYlwYJL2guUjcdk2C2TOnooubRH03U8+QUFKwBuwxHa2XeXpbFgAwZ
5kRVbeBgNuKJqviERpXxMymBgFVuAynms1R32Rz9iop3GcFj2kfMCCBxsZa/JYAP
Lc6DC+8C+rL7om1n1ZzNuKuwA6qU4KoiRtooOWusxOcMlPgyBT77ieyGb6CT3SLx
lV+cxGAMkEpVCQCeuCDltYeUbTMRwFMWs+/+h0RSD0sKqxN5xlpOq5F96vfjNfvY
sR4ZG2CiM5axngG1nC1Bw9PHXuZY1TCfbiHq79bEATzbMEI+8+rBkr7rwVLEv4f3
IcMCn7cw9CD+ZksusK0lUeWPXFN3xhzv2K9wfctt0XIlEQ5hlvUVhm/fW4hyPEYA
XHQVDcJtISErCKWO0SkSxo7lQkXGeO87739JhjWk7gCqFo+Gtop4VaOAPmLF7dj5
4fZsgLyO7xR3tGT3LmJZWYN0qHKFGpoLPmTVPtTmrCCtx4xKIDiaNz2XU22AxGLe
yc0tcsNr73Ra8JJvhYAHAFFn4mmNSg/rdzmg3EGzeg7Zbe7uD1obS0TvP5s2Y4pK
5CAdu6lAZpAZMidGhP9LQAci9UOAqq7maFJNNboZFWU=
`protect END_PROTECTED
