`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0+3nICzYOg/5LgQ5g0dLRcQgBkeq0kscBZFLuUU9LyUlej/b5CXUDf7u0+IvbXQ
TdyQawurfEGqwRRnaFCWVGkMxfrKn0zokfnPYfqmW20c7SrqqjPvzKcvej81jGA1
z2Xt+LZ2wczIabRYOgBKRIpaArDVjkGosnOJPy92x1qcTHLKvozDmmYDUkW1fyES
sn7vNupCz8pEqY5J2GAlwfyxpkqx8kZ0nlseJmwe3QDpDFVbwEQOY07xYnnqy+kA
NC9xAdhz0SR6cQ76JaGsTs7ftRYaHaGAOTxLbfuh5AyQG6uiRUGr9uR+Akw1Tf5V
p8xfKYnalVLWB0Ov1D2ikEiuFwEYYVKLVBpvDGKndKTCajy8aZyJsh6g6fnA3tbW
Kh78Hu7RkVVMdwuY9SVeJLlY/wCj43Cgqw+NNC3HJhLw+IQCf5xPBvPdfGfDuC+m
lwiIpe2UqlG+IQL/nqjHemKC14dZJcxqaoZ4rNoHuZtUVLgnmrImdlwdKDiMARTU
9+KWiLZY1IfTB3sX2p6i6ZfPcoXAit9cNVSAsRJbPUSQTBS4ht7t04WkfDSkw9WK
ya5Oh/uYem9XcIcxqIsTiy1ot+dZjczZwqqxy7S3cDRrTNW8+eKOe3kTdKA2eMSF
sIEzaj9o/CewF2wkMeUoUWdY/M3MMgo2p+JGRDiBcsSRi2U3kSMSywPlfwdrrBwv
bxUn/JNYgQps6o4uVZNJYch2Sb3YxMgQDElaKgxWNkFrnM8vm68oF2nBIrGBMxTW
CHiD3R65a9SYW9YVV3jBXEwnvjP/d6oUwXap8SDJEGlZDqZ47DZ3U8zzVYNaH+Rn
SVQecG0WX7gSvKr81zWPrPLUgRm6+AaP07/Ge8qQvhNEKNSySr8Kpgz7nwvYDi0y
NeAH7mMxDRT09X7amDa3KHLXIjn9eBqiOjo19Ol2d40NPSVTJr9NRL3xZ31dNNgX
9CGBS1CHofot3vKeV+bpxftWcGd2zVHNmqATSlGIxla5f4Nn9tjPSdwF+mmOd5hT
9dB8EhAMWrTYCLUflzmqw2D9MnJo9kNaO4NecVA3YDhk7PEStFsxSoBEvOcAZXnz
BowLR4gGEz7rraq8nxd5XVs21l3Jaysyv8z9ENqaUfoQcvBPSFaL4kKPrdOs19G4
GNxOAfkxdXalmDQaoD2SS2ZPVgTQCBssZLozV2wkwdmIQBv4gTTEoabsrBNfa/JP
2/LXLCC3y9xPLLn3u4n/vas0BUZYPBxgqJ3X43umqfwvl0LXe0D7lvsaUtM0eZxK
wi/ktNObk+F06hcWub3h1zYwR21M/fGqUflVyc0LI5MrvJsb4qPudvc9FG/chuf4
i0P6S5n2P7VrmVOOlaotPohpzjL4N4fmSuD7GsLwGti34L+2T2zpnXfPFJ3TwD6k
I5q9+lX6gXMwH3oD7cy9gBQGS+mWUQE9Chbcj235ZtSNDnD3rkaAOAEoQqq88NZe
/AOcM2ccefKhwmvvszdVBpqX8GRAn5DbrGW8U6a+IcyCECUcFGxS0joUtSOUL8As
EvaaR+pfIwbE+CslGI5b83jQhdfkJWd6usZ1iR1NZCdRbva8l/rAp1CwkKugP5hy
Cw9/+CsjKo1FgakMa7aSw+NAblPPSp0zhMSrHD20HzqnnE0KgArkqtxLUMWZ44PP
9yXy3WG97Gdy2U4YoeC3cVedtdOLzEjUv68/7HtWwNi4vLq4tggydZi25tIEBkL8
8TjbJ9tSlG9li38nUcYAKoaZUxkleZDGXcRXiFBfWL8/eR5x3FkbOVlhfFsLoUwl
iSQk34uvjyHhV569eG5B4FFKKQQEmWBC+FEYhP/XeG2ykWgZfVy1eNk1C9LCRajf
NMzBZ0ShwOFbWMnWWIK5GFvSVK5gQoiKK7wi6vnS+wWEL4brWqrbk1H7I/DLIqQs
p2UkC1T+hO1Arpf1zA8+o5ZJ+Z6AsLRoAX0D0X5DY2lE3dbMm3s+L/iM5uFkLYs7
sCHvEQ9B5RtZuekFkdWGTDEUehOf+OPZ7I0YTW8XAFuF4sVNQ+qzLajwfhThLXVS
TIobFWL9FEmifci+ntm5voG6B+6Y7M2KkdUq7dGc4z9EVgy0iTBhVytgQocT3OPq
q0u8xOXrtqfXUT6AK7vx3L8r6PFfUM0eVZvJEgJ46oYv7tvmZ3IjuZwiWBi9Uml8
/cBObfPrGWeW8At/fgCWGeT1+dBYePKdgoZD1GPI2iPFqQoB6Z1uwmjtCGfrs8FJ
g67YIvJ2+In35mxCVCr4XXC2Zp4dq1G5Zr0xi9BAK8VhHm/ZUhjEOWPZMReVLps7
Z6d5NSXX5BTvdalAyNTKI7E13O8QDGqwyDo4AmalGd/FgRWP1PVVxLAWXTJhc9If
qbQ4CzvkbIA8Efn2WT+DX9bHyCDM9WVyVyU5iKNOi6sOctsto9TSjB8fPTVSz7AR
oiqB0mXHpGCO0vNU+uT/ytntSzVQPcl+XBCTsdZOcZDD+Gk7evtNGOa4MCo5mm+t
Rt7JlsunPcyD1slGxGHb8m8yOyGZmePmBkoTbSuWyvrdssGLAbFk0Hz/Tjx8P0oi
/MpnTU1UOiAMBGg2x2C/iVoJYhlKJWM0SMqW3Sz+7/MRC1EvXyoFDhVihQSPMcub
6KRzWa319BB9oHJYM2eAC+Kpgzq9eN26CHziQWpxCflmNFoXBKSMGpuzZRL76Man
6FAmvAxQwU5QmN/2w6nWuqsCtDLJ4/8ey9KfQj/eN8xUNEFOaKjY85tzs5i6IgUd
5hWgrMrEGiAoOvtfENKoLS/cE9dQH5gEY4eyeXVYFCCry7kfQ7rtT9Rp1T+CBVul
b85rH8cv6pVD0fxlW7H0FWenakuQ/tzgYbXeE91Xuw+wO7fQt6QDGzu0pWGjPCQq
16FmSWshqZHrmciV/6HyLzkrxjM6mldv2DM17+y7OVY8wEt5db4H4Zas1aKtdlIM
93eKVFeBcREDAZfDPyYodn1mlxHMgtvrRRLrJP6rmUiBZNUXo9alLr3kri3EL7jZ
lv5Icoozrtjpc0wwZbM3S4O6l3k+jHtZ9/spffgL3/qRvcqxVh1CPe2fEheVJpDt
Ei3rKXcx2trhmYTv8Doe4sjTMO/E7oowVxsHnLgLjq8O54CKXfuDZhDp3HSohd8x
maDZs9HooHkLnFv/rOos8w7+b9QnjMe7aG1zYpBJ9yA7X4vFkxOscm1aWVM7Gc1p
0UavUqOy9GAD3wbD/NhaMkKSf/UFGZiDhe4my1oetM2kLfVIRT6Wi899XMzVq7SF
7hNL2SeGU1dPmXzikEwJd+eQJS6EvkOM50+cBuBomgnsnlWm8U5tUyKruexOnubc
wgjo1ZrtCMUZrUU+25yaekxw7sLYEe1Bxs+zht8Ip59s3tU/Z8u6GJYtTeQ5sc3w
no9d+/GnST50evCeW62tj7veBR84KZYsy1jBlxZnbLSd/cn8P8LzQdI9bxn3L/z8
8SbQpmAuDlY7wuDMqzyD4pPsg9CHLbVLjro/a6ABRsddy3Y6Jy8buAUgYt07BKel
+HzrpNTlyqgUihYTYoV3aAmitj3BC0RTyBYsEXa1eXkHvH3LI+MDj93QDHOOTxTU
w0vruV7TqJ/1sCTasRF1Zd9ZIyTrG7n2fVP3rY4UZEI2TzOA3F29n33FjiGqPALV
+3Npr+JZWQ3/WEdlgUJZsbUNZEJrpEaxZgt9nBQ6TTpwc5WLZHgvubs1R/5QQa8t
2nUn82uPnzQrOdPRZPGY4dIexvkf+8n2BZyvOW+zzW/bwIHDC7XF8gcakFRO2sqM
WQSmzk3mgcEW7jtM+EmN35olm264aB1VGGVWwSqCkIsGHtWk01rR7ccnLSyeahl6
oSmYuQYfnUc5G4HkW0S9o2Ymcxs3BluVMUbHIbzzZy7QUQKwhCCb2Gx4rWuQD7ni
s2qgZr/Wdu602Vvqvm7kAx7v6sInoqU3KHfut4fJz6PdaEUKMxMrSzc7AAx5T7/4
QZubv7WtB3FzHd9scJvY7jzV9LJ6ALlHuDKJMhKdjxxtuGa82+PFrkx3hrKJ+MB4
/Qxn04Vi1l8E3WwCFCnhyHVPrRh17W4XH2VRolkLW2iUcGQwWKOOQxDH7FgZ9fQE
7ljlEgaD4S+1v6t04434bB9WHYj60NvHy4Pasyc7yueVfovNupDPvy5JmT7wE9nv
4uB5Ei7SHIkcjepmHvuS4QlETXyBlx/ZRnJPXuVtVkFahXQ19j5c7YcEjxc6HRxQ
3EC3f2bpeia8hev/4vJSRht4IfJZXUKtoReEv6lateVKAEXP+dqzNeo+EoN7R6Z/
VQ0k/wUnd6q6t67hKUd2YZj0cp58UV7jYUPy+OeNFDgBRoOpf4DuddaAm3Ve48Ue
1OYjda9yfyTGpkt0Cmdw29l0SjNI3jJfidPvyMFQl89xxgElwMgpkUU4mM8xMAGg
QLw848WhmbMG4DambkTTNv+ec+cx+WM7jiYrWwHLU5WB16zzzx10W3YfuZwNlwcz
cXXUHu3pFvYPxEOXGcqrnosPILsfygBeN4NFvtdew5bYDGqnyxtECCpx+xBZabWA
EZl36O7LPU1ZI1bkbBC22fkD+D43oIZXZq3M78i5FOvQMj1wBwh0XW5x9RVJHQap
H42ul9Lj2FdtKB4N8+lqdeYVnYu1OzwXS1kEBKupGuZk/W6EW0RucHdiKZqv08xr
P233GZwnMvJSTxRS6XU1I9chaCPlBmytZQUipn05l27SXKIYWKGYCZg4ZXQcqji4
AQ/4M730tW/LZvPXCmf70S2uW4XDYYImZNXwCkHpolhf4iT5BUYIW8m1RtcgWoH5
ttr9Mqz2L62ywKAZnEIfuKcOawvfslfNroCrQz2Ub0G2+hdlTp9hdCl5q5wYf3sx
gly2zYALdijSs6yU5u3L9U3UMhSE6QIG7sAeKtvHUEi9U3HDHuYsK/F0G4E/AuQa
oQ4JajAsgV27V2IQ+lfPMfG90PUWtXal6Q+MLrxQKPOVyG6bgx5z9cvg3+QSL5SD
5Mf4Gu0UF8hSuWYCVE+SBry5YUJPnSVyxfgJsQbpnkwJmOsRk++vYAFYY8Jqlw6T
Pz+SkLEUuFkvF9cbXOXp4+AvH/WPuAZe4jzb8NQt30eDT1qp649Ze0K0avPvh/ht
bH0ojmswseRw8Zdg3EGiSzdvjzaipDOrInzOQc5RbrivOq/m/cDpzW8pyanGo9v4
01puwYe7VtZOYaaondDX+VoBhi5uVnKmVsGVXI8OFHzvMz8xR49Cr5azWaUg8pR6
eBBCDT0X9Z5FaTyzA7+aolw9MH6kZm9l5pBnsQOfN+EBiQ3yNCQ9sHIAqVVOxfH1
U859/wi/yNECcC0SfLJ0wmZozapLXCHI8yyU1/XWVG9V75QJQ7SdRVbXrJE6yZiV
wpC85sD+v22JfgJOmaazswc3l2+XOPGTRwJ2DZPIQA9/WcCUogLhvOEJ7Y0TpIgC
uTot+Gnx8OBklJeaOPdjHMaQSLhcExGh+lrkq/NzEKNIoTXUZyaiFf9BkZm3rx6Z
JqWOLngPIGMc9kMhnUPU+5spAaJ5SMcWXhtLUojYnekDe6f6IA9w30U/n4IhlThx
6Mb3SWekrED4imrCttzizXO78MWPW5Y7lK5bNI5Shzs3RU0JffLChcGMJdk8oz7q
whRhT3bqe3Rcql21msG0BgPd2IrR8awjR3woTN6ff6FYXN0A6TBTo071NOSaOMF7
JTizlXUdLu+i07WKNQFhnoQOFnBCFAmS2Cb0EbZj2770mMl+ZthfZBvNdUB1iS7C
h2LUfTldItOW47NvARHOEJTFMBYBcIRevIUt2vfxTDGjBsmB0Jmq6v0081XXcHhw
EhPBmWdVsKtwRd9fd3Ri5P+VAvVUcpLoe5emJA+Yqf5VszrK+E/leq5ZZKxVdF35
IWeKL1yetecib63vnbjNtSePAfwmntB9pJ7A0mRnnVltzhe64T8TO0phBhwakGE0
Kec73TbAH4ns+dpY1cKYUPPSQ76BH0Lkay8LjlsqqVrLF91hyxZG11TR36az3g0O
0WVFhiLPtKJu6kNBURq8sU2fqgcvoDR3Es4hC/4QXkSgLaG4OZdcs3L2bLObU58v
Uiz2vRSL6RTOuEy6aaejTiasTIfTkV0CPGr8g+MkVR355kbd5uurjGzTw2GZLpg3
TBlqcRScHmiK7PnpXrftN9MZ4/FYjkUq/NrMxgymMvgXkXehkIdPMCFvm+jWpDF3
lXdys9wvcW2nCZffpSScZBlyyTmQgIR6aqsP/IB2iOKilVHW9PGXTjRPyjWthX2N
P+UMtQTXmMO+un9TPD1J8rOydl4IcA14m5w8Uv95+YgJCdGIizBA2QYX2ksTmTwi
hYzw/2l66/2A8FEUN8vlI3SGqEs1ubj0AO6YVjlDb7dSxfqqSTejCB2lBY3qeVCe
5/B5GVXnU+cntqf+XfPu8goQW9v93pjGUfM1cWagSUlMxvlYGcsxMjfEUBy0Tg3e
hUqE+X916xtVeLRdJuvXFPnj5eVwVRcngVAYZlBDvhwFjYlfsrb71YtMqIIWlmVe
T3KGclZ88D7cuSgXznRPc1fNDnsewyJOouhyOZIs5U6ik99rugynEUnruZtZkNkc
WgSJqfE8bVgjn2kUUSDosQfWNatttkCfzVWDf/7A+0/1l5bRWRp9g40QFm8IF5za
bg/CnoQ3TP2GFVccy8/GFcwE8a3JWtFO6kM4VpbyfoyRK0Ye6n/awLXu8Y0Xgmw6
gRyEOFZlFHQGJVK6Z2xwPgDEY2yIjOCiP4HZMtwWY1P9aFH/qieB04jXKOP/w+4/
H8UxQWMaAAk3f0UQYgGl0aqahXTuLwxo8r26zBqbepxL/xAF+JO3DNDkxzQWdT4g
+zyIjka4w8bRKSPDs8OyxTzxs9R5qgHC1gUnw/tovqbkIbauENM111IneQJOdIQG
IBXNqtAhHtWZJpV2xA7Q3bZI9p2UNIk1CALea+liiFbt2Nj5rm0gcmOVNptnjuBJ
LXQqIl+RSR8SS30Y4J+HC68WeO76JwJ4fjaZ30Y6T87PYxEje37tGxEvFy+oXS0J
zY4eZj43eJ619oBNBtaixBEh6/QCafAjStHMLXbuJHE/aF4tzjjHJuiwySLl+nZg
p7WlYiy089BQ7cxR7vlYW0+LjkchY0bfTCA5wrdHnnUfeGGWn2wcSkR7+PbUrMXS
gT9tgeUS7dRPCX0vhc1zQxhAd8HiWliXJFHyK6iSnVLPkooUk6tDNMDMmqJd4tnh
cJ3ac2+OC7PYNfDrzJahbwWUEK+yecLgMCYGHDFgxBVooGZbEyi7fF1cbaHsvKMq
bFR+dKhuSeuYTcYiVxonibvVBgFlYkcEDL+YvTIt3YEUqH7lVcP8JghLEiB+4UZ2
jzhQNAgvNga3MrQ135/nRCOfRsWyYSOdTfzoy6Psuu0b8Vpw9HWvKREyKi+u5WKp
D1FPGQup+b+ScRKhATewRFEPQ7RPkBSmb3ODWG6MRLYFshwl1RJBNEgecSR6mR5f
5K01H/INZES0FEsE96LHVNE/uYAFzsLDSE5WmN5zqdgpS0hamrxo1s2AbXnwRSNL
NTlYMREdWxn1hJ4wUlUgoSd3Nh2DDONn695BEPEJPueSnqWVvu8wyNeYyQPU0dGA
H3w04NpJBKyn+hgBOwh4ZGXHMweolM+0dC81P4Bn9h63hErCVCVjN6NoYaoC0Eyr
NSrK53ZkoeiEnkeSCjrH4fF/scMKq5tR+NaAZ4uQsKnt3Gxp4D4U1rycSaNEoqbx
rzScn/9xQmk/z5YcOoKJn6d1tJzfkIDbEM5O8F+u0kugWhMDlZFojD7S6PnCyGeK
rtTFt+uExMqxBf0LyV83B36QUomFvhyxPaqGSerKhSHECiNZ55/CgS460Hw5nISJ
KBp7vikNMsbAvvyzUM+9lZtBSgneosE8nhD+g2GUAopMxPWBPsvZQjXqYHor6G4f
d2hr+Yz8L+eVruoKtM+Vbep71+JqkGcIgMGsO8DqYWsJUOku9wPLAM56JHM9JpgL
l0hFjOQ42QnIxHpKnXAv1Tg1SEd4VtNMbLCyUrj95dNuHKnhTqAhYeCLgkTd2Dpv
VaWGKaWtBgCYKD33VbK99V53m9d/e96QehIZvqiZgbZ525kWCU/QlK1nYnmlJI+9
0ZdwJkEf9iubkyG76F7D5xGlvFx+zDycn5ZqepsNXTfpV1SJdCqocp3XCYzmPmnB
pO9oSIZ/wMyYb8Zq3ZGlJvY0YAcs6tg6B3XW2hBIgvqFlOhfVNDgI01i12PtiYRr
aLtt7d/4VN9LwH7dJpicp8tcKmRwxH5Dud0N+gp6RLorzBCCY2ef896OLF1DtVZY
hG2LPhBe0Yypb4t2oy2HLP0kYP5yiAaZYj1Iz6IgMtDCu8rjxbtIWVii/Kc5ZYYB
kIQksURno/7Q3GixDsgfztOma0Wj6/OOOjMFFDGyb93hQ8U22Zh66sNtg/3B0PHR
1iBWPbf48GZ3Xm/48jper3L48l2HnoJ7T6Kq9TrPW8fzKAFcmAV1OaC22DixIMVW
j19aLxFun9hzhtxdpjIaU/kb3131oY0w6t27BM8NSHKhiI6L3YBCOpBTkZNTwPjX
deODh9qs5GA8vMAWsGbxtk53B6tAq3g4OgWEPQJt/4inqZI4/3p3JNjRO5o6vS71
v+PkJNdhaU7b7sMD/y7y3Efym8ih0wPH3wznsu33XUVbnu5c5/GZa57TpyJLYyPg
BnHBKYMdCl73WM1DzQ+DjQaGHwjTMDJAufwi9Ri49oOTa2SoxeaBJgAdWLzyHJPI
FsTvefQwQ9+p6Lf42Ucwxhu+azc4PnL1syYScuJsVDJOdgDFPhGy71ZjEJuim5FD
FYrXIA1uUcJ6hh/dJG3rewSQIcaG9AuDIAtJMUCHHk3IeXaQvvTYj6EuQzm8zHDZ
r/+HWX/NJafJqLUMSLVDTXsLiE2gs+R8T13ViWkCd1jKFx/AP2EIpmEW++2okCvP
f1vHHOJhJgFMmue62XV9E/mLasKv2xtAex0g+sST4hhorpzT2qAedKA4g/07bOHu
XNhhj1a96yXl7Q9IyV3Ah2m/An6lUzx/vmGuY2kPzwG85J6pwqVdBveIdPJJ4hKd
f149RJlSUQhV834WlQ4ztDpCNvotB7k5lEOTg1JJEIPtAkW1Vv/1xNoFg//QTR0r
qRAQ+lu7jAuJoaDQYhJCngGBkK/0SFnUZG2vAoHmYTkQprJ7GRcoYhNf0uC0eYOZ
gUzj6/uP4sxCYBzarfssYEU1Qk1/0a9IFaG5i6UTwPa6yDcjHVftAnxebXo+YY2d
18wl4R4CCGXibYcYcQPw5wBppY06JZjQCkrCS2E94ZPukYZy3l9K4viM9Hmo9eyy
hBMMy7QDuWL8vGkgyvm+HXmTdhX18Zg0fSQj932Wk1ZhOHzI9XnyWH3NAvSCHPhn
U34Cu/RK6rF89m02KWC7R2vaBh7ZaBgqYEJFXy6rUV7qHp1Qf5K5CZ2EZry/G62f
p8BHYsUvFq6SPRClnJDUGyJ7rzdzzYtfuKK6pg0mIrjnxsudos4R8wn/xu1udkSN
Qt4YLiYINzxqiuAUU8GXaiV9JoZ8zlpqkvyy/9k+KHMS8vJP1oLGwr7Xt2dcmEF0
NIWqLTcJjfeza8dWG99blBNOGiXwS5X3Qkvbc2RfD/QSFWNATSj/Jm7A42fJQei2
/0jFv7ikpbzMm9VQJ7WN1umZ8E8GvyMnxUveAA0B3TbRSdTM2vAt4pon9zkr7onD
+ha1+rOxJkdeA96CURDN0J0uids7KkZ+UkEJV+oql87GSOo+D2osDQJYgzkfAlLy
rVPh8S8rDE6AEk6hmXwhvucuyEfObv+GdsFnb9zXshN4WLMpyrX/Smr10XS+tmaC
hCPBEOTyp/uTaSxRc4bEPRMFfNI+pLSGOu4RyU+gnJBZ59eKc4runjKR8sWmQasx
YiuoabvPCWc31tc3Nq0NKMuRkB/JxO2LWZZeL0OxnlGYG7BUnst1DdYYut5M0wn2
kU8IQjvJtmSQtE0JoOrNllmX5bgegCp3TytLWOJIjsx14Z52D58BLdZivjC68yKe
N5SZ4C/5Uu/L3yAHvPqzsJee2+gZvOqKFkAH/VyM/wUhPOneqMMBg3lH9I02mQoJ
qJxEsc1S8Wjnz2yH+ae09T72TF32L0bJlK+nNeuMBYHiURqwkzoymZwW6Okqj+yj
y6O247wBVhGtW0S6WGs8S8ZorzUYWAPvkIlHnBxhGjDOnYoc+WNkDNaznkKFHq1T
0nq6HG9sY4OA2/JaY5kd+qUOgTJuETNwKk2mEG0f4Ww4+ulqqLrvboPT9RLXldAq
FdZ+c/kfS5+DXxu951aMRbQE3JKNGbfKHFD1EDJnHSnFjIVR6H2VPQrVKupIR7oS
xntalQGyYSOGBF2QDfqREYC/gwEqk+sCwjwXx4ofD4SgsauWhrCf77Q8MZcveUaJ
Gh0PLNDPtPaqkBad76Oy1DHPpm+D9JgK9QYprTK69zU=
`protect END_PROTECTED
