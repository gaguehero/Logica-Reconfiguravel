`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwa2KawmOpbf9kUrgEx/uAq5RZG2fa5yx44jAXwOIfINb3XhoeiuethQP2PzghNI
+TecXwpbt3NAuxBECN1E/NCuaEZu4/uX9p4Aq15AyOxXUwi2lV+s6MCg2dbKRsUF
tgd8mOao9QQAyIjgnEaMVdHL/N+xVYEKX+68Izqrx9q97pVxtL2ZX4XbpOwOLRpi
W2rd1XPOkRmS4sgK2BxpaBYnvicfzXDvcEjNcRXoOgtyflORNuLdjyNEuK9fQtB7
we5KgkkfO5GrmY5wc5ThdhmNK0bAQnU2VP6EXzDdkUCES9KonDZiQqKSO4mJZLdJ
hJUTUNGaZei/dKY+tZrFQDh2M4XlTUZAL0vP4r9PK1UQSlEAhTwwAKlGKQh8JQYX
zUh9sh2G7qujoN14tYvVk9IiVSkUYeAchHJWadkiM5c8//pE+qJvPKG8/0IQTCXS
SZKwtoyozuxKOasbyAR8iU/fdyUabmKDmsPDl+gSCzReKG/2ZRonCrrq28rKS1sL
GWVvugxepOi1OqJdH5S9h39a174J90DDKtgDZfpMGf9G++ntyh3pgpCcVVom+Sgk
HmIgI36rcCB6AulHEEI2RSrQFcrXPKGfc/tjWsnPNq4KSgTzrXyxEMZmVpwq4mPw
KNk1VtbQXAB/n14ZcD0uueqsSSlPq4WTYGmlEbWPGp12ZKln6ilSy89KEAiODiAj
Fikp6P+SS2gsGyFeNleM2ZhX+EGGT2K44D7rjg/3AoqYTzwwjf0pjyijb1E/S4J+
4lwiER3hPEbeHn/wKsxYh3RX3s4NxfYwW6UmqMpcM8cN1HFsV6JL/c/GY4uLGoC7
snBsNUZWpPUB2OGNbv+ZlweWxK++EEUL3g93Avb4dhhaXOy7tTcJm6uMHXblCyeF
aZoF59C3xSZG+9FhoaGh+wgd4eRamueZwiD6g7o/SoTDPCXgbThxDgpqHbMtAULA
KQSoGhlMusP/TztV6Yk8kkRPyQHoWY1lHoQZq1ZMpV5JHLmLhX7v5cO4js5rfiWQ
kBztw/iWPz0WbFlKrrXOktRZF2X7BReGDBjACab2fTKFZ/iwjK0+rvCtZZxlOOoe
6X/T6YNUdz9DhVSg4KM13/NBW/C4z0jQTgmWaF/t4LDCczWShW2z1bfIPQEJBGm/
Y0vrRlBoqLQ0subTVFZMEIYiGYnfyyf0JZ42N1rAzULHM88KeMD3TratwF9W5QZ5
OewFeZI+O+nyO0SgIEWw4s9+0iW/3X0yawjcCKiOlPFMCKS+ttsvWI1V/SZQ2cMi
j5H5JRh90fFrCaQnCBprcJmuNUPuJImvJFe7xywM8SPMNYqRC6OwIMEujowjVwGU
zCDPMtDxlxZt7sJU8kdK6nFU4xRaFXHKxwbpQ/Dbc+vtV2YRVghVOFESrFzrqiKT
tEZFcRueRYX7FvefE96VgTf+8NUUuTz8b2lfN7fwvTom0yKIxyKygGBZ1OLWhFAV
cXsT9a0aKf1OhHWx5DY9Qv9w8nzHhb5WLDkQLAOuJInm3ctZzF9Yx2txtxOncVoj
9A6cqpP6PV9qbHsDpOo0/O/qcpMuwgJ1xnPHxCw+WjJ9QweIt3zPIWVu7uKZAwQl
YiHfAZ5tScqrrus9DNIeOdHhFShV/S2N7hds6UjTh/tupGGMD++XRd/3nWx55bUb
ejl+2Dse66YoZCYQ3qi873D76qTMb5mobdw4QVKNfKBh+WX89qSKc72V9ke8mu9k
Ytyy0MibYedtMmrZfz/7PlmFGG0EaL211xxEJsix9stikIW0e+571H4mwDDnsK4D
C0+37QATSsD9b/SJP5LE3CfZ/EqD0swM83SvYPOw77AElx0jVrHT1ibxP0siCQJT
/xTuiZiEfBLE+x1LTZuTzeTX62LqE37eqx+7l3L8RSf9PoRVCzHuOjkzWqQ3tOlN
XcRqQbKd0xs6MOowH2Sk5sV40gbXsObLTHVcKFsEIWT+4jqgRPNdqBTA410YSrkS
m6rwZiuO0uLC6xndVEkPR67dE5y17PmGSa78KnB7JHLGonnFDKeC7d8TBZf24o75
YpVIDzmvBb9E+viYj/rTa4QYBhvJEcocwEPWXjMT54+BfWWc6AUJPhWG4vw+IpMm
btzdYiauBl3wXyLvrF381gDP7LAotg8VL+iWL7jZaiqqhRc2ByhCnY9obtegevEK
WKGHomUg0n1uRjS6Orzut5nyd4rlNpPW4utOH77m9FHFDExrvartquXb5WvWVbSx
ZjKj+x+oe0IAMff/WypQ0LusTOHTIFZ1B3DtHj/INP0OUmW4WdFqVcmfFsTKWbp1
2NJ1SafCOPvey3PzXKty3Yiy61tWZd3Y2kLv8eLd4jPBmYJNlnJt9sKY2h2Me4xP
q1hSMe94WhdWQvLdWFMO0zGCe3PLeO/K2EBUY1nLqo29/4QuMHrAd5AYp/w7K7z5
EVxDqDhSjulZ/1FDPBgiGQ4V4dDwzZfm6Xs5X44ek8u3fk5F5ulqFqEireARxwfB
QrtkFM5GF/XHeOTEP8jKfIUx2u8faNGndetJCueSD/vIMx/CvZC9wYgpwObu1iHw
oV5eQM9vEUxtTOdgFVEUlCay2yf5JKmPRjDUPwWmX3geIc/hSVvHb2IZKPhd6ems
ZAY9+GRb+LzDLKTWrOXgbm7KB0MSsHT/gsO8hDhbpwDPEfOC6V5cK+0SYeHe8bLV
+XZAiSgutRB4ukjyniKYS0E8vSxKwPpKMU86uRrg6+y3X00WWvLB8aTruwOS9YPe
ERr0//BjC8mTfafqswWUFsqqbuynze1F+Th4Ai0ZcOZML9ndqn3R06BejtKgqZU3
MbjvB5JozcoWZR8Zoz75WTvtnzPifQS+Jz1pfslR6HzXIei7RBGJ6J5wIwLsa2S+
x4640pYaPscGNtmaqOaFw78kis9Q9MIcla5sbEhibuoj0KVT3CKqSE+pfwFcJ/IJ
QscMUNVzWMJMBbeNqBP3CXbNWY7KVW01WRwiU8Z6dIPU78nZz5tOtTXlC2NgwQAV
rCGA+OTsgnf1qTe/qTSROfZtIk+sNDTRGmWyhanee4j04Ij9fhuDFedhAs/RKsLt
nYqQkefzeGt+nv0Pm0NfLGyY5n8CvNr+pVL8mXhbSKCWafSqI0Ak+jWX5w5COGrW
XC/LTqq2LsZBzi8ZbQ7rvKNP8LJrAUUP1E+bNjpMihYnWxof8qP048BSVDptCl0C
+wttZR+1qkh3WTO9eOrDRCvQxKd0hznGcpuhbLuOM9qEd+YMmC7GUDyiqUUliouD
LKv8vc7/RypvMWJ7nbRKDsVoJSApzN6bLGpX7fq0dMtRz/4WMfl8TF7xthBYumxo
Pc+/TApHwKu6zzpFtNqWqh8BSqFmrC6mjkxbL9hD794aVWxloquwp+WeQsYFr/R5
fEWd3Y5zAQ9XthlvY98GoFOpmm/BmEdqRXt9us125crJIM7Nvqw8cR1ntPnEAlLf
YFGJMNCGs1eKZ2+1MzWwS9qn3CCN7VWLdJGz8UbX6TTOdOWjAZRiesZA2gkcUQvX
mBoLMmsaV5x7SB1M5zLs77ABkGrHhR4eGkNTAHSrtgW/wJoruKp608B4Jmb+92so
W7oU7inzVHC4/cAh/useVCMpNnkErhZ6QT1qjOKzQfNbuv0SUSQrlG57IOzw95Yy
bll21BoY5+CND3N0+iVs7FIZuf301/cE9shuLoYjDj4Q3CTgIhIj01D7iFsvvIwF
ufcld/JpUK/+s3xcoqRQC97UXdFOBpEcatIuQIEUpaI+L5U4f6zlncfu+zpOI33v
IpRm4qEYThuKWiMvmLLQxsGDLVPVKcdNsFet1XDki3L6BYwtQOOQeB8MO+Jg93Y0
SPj1b4J9P4CZaUZ4S0CFCUKS+UWtD4ubPRBKpc0joEqIpOi1zjZCks6vC4DHYmME
kJFy3bcGVlwq8pc9T9FVXh3pqwWKyu43U16vRsRLEDif4R0IhBMmB4EUe6ttWMAj
a0fiVFbyfMgMU6ENr2Qz97ZS6FFeCdjg/d6EeMqfkcU1rmM/P9ZRQilK1G2MXAWv
qbnjN+mmYZZM35E2B7xfSpf/oKwNrgkxYFEp2ISou2GuzjXUYyvs2BMRBvMqdCqQ
hMIGfEYeA8H+NLWsXEHaP9pPJgT74eX/RFtNCjaYvl0wq+OXOO90QJky+0TXPh62
rWWkbX2eMzk5SqbMEHmwo80u8kZ0YNDrmGw6nGDi8BwshOaKntk0w9oTqN4swpGf
SQwrGKG0u0RO35jlHA5jeACm/fnAKcH8nYsw8zSw1gtG22zBqMk29Xo6BrhKfDpS
PqkmQ+KA1hXcxDJOXI78Ns60WCo3vsbj21vLGKpu0mran/eypBIB5SlTBkvvXvQs
lKbc+8R8yNJZ2unL24NacfjA85HR4Ohdkwmd/0Vkk3VZdhyOicYEEjItkGbcyEA5
Ny0M3+LZWIpiIFl5NkEBCRfqd1UY5L8HjY+L3lJjjWxeq+0/qaWTB+nqeqdrnewv
V7nq/YtgReGcDGlKBtPCcMZnjiSiFVariXid7vIkgmPLkD+21mqSsLLePGGJhAEk
saBs6A9oE78Ql+oK4BSF4ZPzZ4rBs/fBTd+crI8KjDkA+51OkCh/r1KPjrU3K9lf
fox53USHOIn8+qoqPA4MCqjGs6+QaBYmSZc8NaVejzKdsXMbAcantVzyshTvwcTz
5B7HcIW8VkCk70mxvRhVT8covVOIxcebeWbiEDktidpqVFnCv0fgrrXx7zv1NIKP
GVWkX2qic8vzmUOWnCoqsU+n6yMAOplJ2/+XmBYwtPN7Uj683J+iR1nisPgmuPXt
NXiqs+099VIjgAh2H+sabqnlxhOqYYY4RQHoMqr8QG/dlUJ4S4wm7dKh7+sdNchd
EqlNxQ/S51hXPAuGZHg2KVCUT2OelbnuYUyIjo80G8EsaAIDNmbCK6kZClHfEQtd
BUFICDUi7+RbxqpG3WEJ+8YR27UHpoFBUSa4kdSBBvCAT303xvr0AmSZCjb22XKz
9dThUwAUcpQuHAgI3YjQR8viGLPzOHeiOyzjk4Lyl/gj7DyX/Yz+JHw3ljHfqY47
NOnE52HHseQwN1vDP6216VhPy07XfBDz8m9x4svnLGXLQRzqvdv7EOZsF5WJ9/z5
sVdCPxZsEv3zz8pdmKrp3VBeV/TgnEjafzD95zeLo3YQbLs8CnjCh5Y+0euJItVM
iqvU+GY7mMyDQwdcqVHEmGScazL0LbF/NGD0CIJWSaCe++ZIjDJXESKE7SJ6fCpG
0Dd70s+pCPvOKv2E9ywxOdW8AcGTGikdXV2sRtlL2eOyq4PJiDMtFGfyvYt51/x3
QOf7GvT0yOCTjldP4bP/Brn5bYtIt5Jjq8k+shXBKOepMVwaXO5nfLWp9iWohzZ3
/bEIxenY+pRwAPgb8Q6mqU5fG1lzaRBK9XFtY78VYJ3+5CP+ri8PTjZRmBx9mE7t
sx8SHZsWo66EwLAjlfNb33jiChxAg4M4z2PhSx4RsEkxRPrFbSg9B9Igz+WlHP1y
VDqtVUKGSgZECFrLajIa4nPp8qV4mKigM6qP8qBkq2D+BphnoM+mZR1sF7XDchX5
ZevyI3UNkCCnZ50LeqbID/knIe9CIpJh8ZZl6w8RncW/lMQavoU9Tqa72bevqB4W
zjBsqIf09WIiN1rtUrLc0io9oUrEV9VlLc7gxuYmprMH9mZAUGz3puBfkg2kx0cd
Jt66PPnG/irN8s6Rjbx343laNbAFVoBiw7sEnjb08q0R9HsWkDilVqkOjPGeMwco
/p7mAIwZpAb5SYQDSD9h24BM7hMPeZkkbgWnfkVTElFtEjkfnkWoMuRMInR+U4s5
fcMhIfg41TkTXB0YHsXuu8eX/0y8gszY0avG9F06dVgTAbP7Qq1SCGwlDYbtHoGE
o65/ZWNW+SUawiw5KUITsQtM2G0c/s93Xco2ygbwJYEB7G+f5jyb4Gn1sSOBDFK7
D/gBVN3WzE2FRfI840to43H/92BAytByfi2Qowx9lWwxb7O3GJaUEES8AdIm2ukF
QAi2DFV9NVa8CzmvIt5hRK/Gx3sx3HyyAlAjp++zRqaEcPs2lZDu1TU5zg0GZVB0
3tvsnfHaJJ1Hd73bd11IF8D79lmeKrKv6e+AGe72vyZetWX/mVQrJLXIZ/Rx1Msu
7COq7meWgiVNMMfh0BvUafvf+XiRCX02h0QAP/is2C+lFViS/3Jg7sEBkAaH9zKV
rhxu8/U7dtb1lAhcgsbyM5W69yDS1G5K0bCmwKT2Cg1FFxsSD6tTZJYfaiyfdQV9
bPzFES6+0q1Pcwo72OKIl1AlHNyDF1IerZ1r4rEWEuh07hqvfHu94GMgi2nkgXDE
SrsKWkAVgPdFlBJMtMwylGjW+FZGH3nSSFG2O1mLzgYoBIL5U6umY5YJ9IdRNRdG
bVIoTAvY23pOIB4IfOi31KAkqHHpQ153jObHIAEF/hveiLRJ+0eX3n0iTivuRsQD
EPe7KI0Uj39IHgkI43wVUmuRGIeoink5UIxnSsdE2zzfcijXnBuIORa3kvO4f/O0
KobQX4wJ2QUAa3xlKHYBfsBzAy0KSRXfvzEv+CVsn1HfAm6nL4Hzl2+lYQbUh7Ef
AnHOxIsg6E7WJE4meJlG8FAO3CDtYNF/kwuSR1Lzt/IQiJ2Czb8b/k8klKnVmVZW
gLp6HkvnNbj9rC3y7GWuQD99mn3p5sps1YzdAWFXOYtBggop9cf7vyOpYYBK4x0W
mXhZQ+hGWcGowxiY52KISz1oBHsuLU69aeJK+InUNKMfJ09buu4Ei4c0E1FB1tqR
phQllO41knbm1DLvZ8/fhqXiKZXk/7zBMbiR5uRPB5m90irDm05UGqLBh9sxEw7w
JdKJqUw7/IEWRgcuKN9VwBskVYK54ums+gziglqayZp3HpOnmBXs4CwyB6JyUy6A
IK5RN5h2BO1whX0jbFwIPBe1l/Fs7c0MX5uZsVSDyTKEZKBeFA1kdd3f2LotAV/z
/KyxWPavnZ8nuAIgcN78cYFJUX3Wy3lW+EEI1gir/kbiYvkg+nldyhI/s4+C5YgU
5MWLTDG1gzaoeuEPJmg3J99NqP39Jcb+uLe2NW5OD7fl5ctNRqCckrbtXnxdkM4S
Ek7buiVuNgIyiZFUYlA5t/mqUMZEwIqxxpDeTuSfjxXloPt3rqwX5MjJc9cQ0TOR
vu2/ZpEW90SV6244HB4FaF+VYQIlosL9deFlLvB2E94tBJNELnn1HNuirF7+HmYD
OTh2VuHssFCGSL2TJ26GyUnS2m8ufPYCH3DqX1WevD/ldX0Uw15dD0uqb2FksbA9
A5FT7xDZiedYzm2OJsLcJq9ohxSNzh1MNGCCYLlv9ZRgH2SyCr4++reHXryMW6zS
9qWjxUOOd8wBW98R9vgplSyokGTC92IXbQoFLHJO3Q298WChSbx5xFQNWI2pgOhg
D1k0OLAYHQ0+SrHrJG55YO5AuWvOLIu00F6LcWoXBk2Ko/AD7/vwjB6dxl2fpN7I
lICexTAtS2XbVOjqH7oj02uTT7wX3pujYeeSvNdHTsUZpM2EtSv8+vQkz+SnNoCD
r3fErmfCmLmVlZW4lrRLZtW3iis1YSiTSTQc74rgRUJLQTrv3MPraUP/YKX+sMYo
Bx/nGat5eEdKy3mwLzUzXZVAu4Aq9q0pifVnbYK03o+RF9/uC9c9v2aeK6aXDoFG
`protect END_PROTECTED
