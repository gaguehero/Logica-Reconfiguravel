`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipBZFUo7qgVs11Wv7FDMU7KAAFGYHH1YEzdWRQVXc+0/2ts4g4vOardt7RzLAAZV
IYAYxnWHh4LsgUFasbKK4ifhtuWnsRLQyhGDfJTz8eHLoK7mTRnmBb6S68SyzIAk
1KlimMrjSkLuQsPrd/F66qRZKNXOvO/oTM1vu5WR+PfpD6xPqBSVUx6dQuyoFi39
WJxVDHdf1A2upZtNnxVAuKiKKoT2bpehaWYKNPt819wqkoEhTcibMS3NYyElbQvM
G12ng8lXQKD43y8Z71vG5V8Z4+N6TuwiuDjDo44Iq4g4GToSj4KAKmT8d6wjrF2s
jQ6kchhmmKVaOYHyWVr7nOtIp2nq+tAOBW4jT1AaLhbmVUGx2r2eqpkptolXksmI
QP9UPUCSYHB+7SmlNVKfK3pmdDd+HshQfhyrV98zzeo485tKx/Wyw3ThwK6VeUMF
8nD4bX4aCy/oQn3kQTrResLjYqHKAiKNBTbr18eneSRWbJCy35CQrvOdq8kqb1x9
EZQi0IMzu0p7MY0vmiOxD0Rzkfym1VUNje7GIZkpw7tZ+hiFj4jwOAnfz/IHMYK6
LSWgqBEJKdCF3l1uEBJ3bn3tdePMmSzTWMXhc6wCEa6F3M+kGpb5OjtSv+/xM9vH
wIKyAiQnBbOGnTpmVcVfBpdV7E0S1MptXxcrp/iSu+Cdsktbx8z42ZJ5gYz2A0S5
psxwr11BaHRtXHupwal3BMNNxcpVRvoKP1x5bWqjAv6Mr11s9dtZMvh1RGzmKpCj
uQ6OajPeP2EsgzpGGgdsgCZNVBC7GgvmZv6pm89wZ2tPJqDqN3+KsndUUEbMWjyF
l+V9gk2NnblSDpkeHlpGxnm6UzUpO/XItvzoISS6F0oh9rFrMOaDrDZj9X0QarGj
f3dhapocEDjsaTrqOHSEgJZGBj/CvTqqP83jTj4Z/hMumSK4ea0zTqeswirEHzaz
JgwN8pkJMx/dvqc6iQ5r/bOPhKFUjLTO1udNDQjVULc4Yc3uR62/URFjR8zoHDZ0
BaPxO2wIahZz6X0mYCtNVp95CHU7TlGwADFvJiFKQdtzYZJa4zhNKM8NtBMbbrfV
iTKM0g5VzujygR8FX+3h4rTm5aZ+ZWicjttUKT58yt8bUwKdU1k7pyBEzTpJASgP
3EvLOpkTs+7U/jIcDHdVGd0CReED8JoThV/QeDQi2UffAMJg9iK65l8mcfc/HsDs
pBnsfl/OnTRl4iPNEW2lLKilKs0G1X7PD9p2PZAMMm7ctPc/rcK68oY/0ekwTRIO
VHJj0LTsf32C9a7JUCSIYb/CEHsd4uHGu1vThueFhU+vj7rtoFn3xoUOdKh2OZn2
C+dH/5RYLlRrmqwoxqZo9XPZQBWuwqAz+iIswzWoWCULUIMOwm6DE44AIWb5lLnC
19WUzlTFbH+jeLDiroiuhZWjCA2+blOD3OYsuvJj7MlIc6wr3tkCVTMAeb+Esfvp
HcYlpRqqxEzKDTnLM4XzplEqYo4zxkWj9xZNKVHI/wSmCLvsTWvm6DRI2xp1IbMm
5KrQ+xuH5vmc3Cy7AQFskHx80znUU5+MBVC7C3HXCkqqzxDK6fP2xwE6p4s6I2SI
LVETu+biOVXG5X7xx/7fv+c1yxwuPvTt9oDTbA2YNdrETGYoPhXyDAvH21ObANqV
8qRoh8sGRdeBMBU4q6eFHlHnubnoC2gWOTOVoFQ3vgqtAtKUsaqwOpQZ3uX1gETl
j7h6JjeoHrfNCmkARN407MuIgPpIGNBD31+GZCG6RSdQq25lg53h5nN6ZJONpRgk
9uZzU9ffP5/vxabGZ3KEAtuj38R9hVZXR9c24ZyVshnIusyT6TIsq2G8bUh5Bf5H
Z8C26rXpNGucSO/6wuvha6uZnBCLq8eOgle730q0xRwXgFM5W11+mnpimCHDEUQH
vpkldoQ6qyQ+dFPFWity0NhRZMTDZi7qwaaDNDt/27wzQ4+FgogeYKi3/gJUlcsP
ZZt/K1OsQ5FIWV4jZWu2R5VMYRkxZVksei8xSfCvwQQ0rkrbJv5tgCCdTf9dL7Xk
RzM2n1dkrWQTV/JV/iD6buUOs7VQ+ZPXQ8WKgbvdR6YkD3RgaZSmuxpwYbt1FIwK
fHRH8trPxJxPk5Air6me7Y27xidyQrc7OE7JhlD3R4vK3oGSuYtKUhRwPMTP+43c
UQRjsXrC/38Hve/ZkH0ZcrFDaIQjkVf/CQXbRsp6IG6nkdaC5hk2jUZDUWErf7r8
fD5M6OFMotLsVUEx105Ueljwm2/hQGyxbvcoHkIdXt5/lph7lWUM33SdIe+zT70T
7Gxwpmp0Kk/FbHeDwbeQhV91FCTlU8bunt81lz3t2Qkj6U4rJ0Y8965GE/WGvO7O
vAiyYveUcayyZ82EXvxVituLhsCpk44iYL0dEaf864f0WWjuZylxaKEKm8y1JRsk
u0wyrd/D0MRm6wJ1H48W1AT0kA0RQKlLPLPGgskO5uccatc6l83r7ptoa72p/mN5
Q8a4wWqByPFb+2hny66QHqMXUrnDve2yHqxE607LKd9Rdc6P2EKySrMsy1CwxEnS
KSK7+sknTKyB6OVRYGkUw0PgkqEMq0qYiXT5ObKJSGjRde7aWKAYmoje9Xo+nyuR
gUUTcZU9NT8XHqRrNA8QvlYejbkutkIbaBlr2WmieuuvkVRyvCbgK/kQ9dkMBZs4
7QIo5EoSWW92uT6tl4DctGOkuoHNRd+/tTPPfY6I8k0qP4eTzEdlP9IsLMCYVWDg
tQhjSRUGcqVkZR8FX2NVUhBCIPYb9irxvpSe/XbLKOXDNA1M5QjfvuHT6/al3r+8
GJtcdR30uryteDq4bktuV5Yp0mbJUSGdo6+OwemkztzWpp5UFk8+hYfZhZgZeyHO
LvWZPe1Q7RqpVc8vsDiSN3xEE2HuLRHXzjeT95AK6wVzx5+znM7nC/rrUpaW4FdZ
zfS9vK22Yxc0xmwMmJ1Nmvj5bsBxc3ISZAIi5ysVuQcgkbkqAhByJC4NbUrgeKNF
fo3V9QhHLnp3nmDtNr/y/h+b7ceL0M1UTCXzzNEupq+HogZgTWvgk6IEetMsCR8P
gDCwKVuAGdnblbYQx1KDx0LKe9qwiHI8RU20dj0lEOxM8unWkMluhojgZZ7G+au3
lxiqE+n/+g0by/FrVkfyQ3aqKsDC4YY++jbvT1HkM36MVbhb2NtQkfZobG4ULB1K
s5LO+uSF+hN7E0ez5bVoZ+TeVfd0eYBV/jdQ4wfEuPn/iq0M0YtZEC2nePN74TOz
TUhJH0T46yNpo7Mr61ef0I8uBsC+1ue8yMvJJHomGUlTd7402D8ulmYO6lZyOVy3
S1GpgiOo9uE6sLvGqAVFqWb1G35E1R9KxZlq2i/Xd2KWRhbcitNsYU4MkYcDy2+H
9uxAGd+0+FXxt1al8RhQ/i9bdXi063x22+3jjvxTycfjgXzAldfJJJ2+rWhg3xRb
axYQ07M8dvZEvKrC3fQ9WcIxaxaoRRRI9VL3mFuMOBviVIe+elNbe9i+29sK9v+k
zQDYR89TfD2TThRSbubxeocwYBvVDrkoAPwfDBscQ6HtgruDSXeL+QXzkv6lbOM/
N38aQsOeVV25ENEnGimYyadQPgYE+AC/qu64/db5Aq9t1WrVIvhy9OrN02n/lTnF
eQzcR7gXlLQVe/UO62cz5r4p+7QRN5Z33/kOOclAhUJzWYvAu292n4muRcVDMWLI
TpMsvVq2vyplZ3vZh5MNkySzV1SRe4qZZVwXrTjsCQUTJGU3e/KNnwgeK+0gh8mH
jpl8FNKv7ZyX2qhRS8txtOqd3T5/dDa50JaR898TZMCDxdBnJXAGWpl8zKX+mxW6
RwhYCQ9SkJdb4/te9ceKJJlgSC/GjQFcAoDefjCn6nOS/+jOjIRQjoZ6vzjG1NEY
BCiB7f44pwL8njLZp3H5kbyl1yHHvrZ7cA/cwUkly/o8M74C+Tu7JWaOYw5Xw5Dj
IuqfRbgi/BvmnxJCKuxhru4ExmXUONYY04mW49UzPg1i8da7eBjNqZDgWkd2YApV
CJy/c1oRCgcB3SLkbjmY43kc9X4rglVQpzrPbSfTZpdI1p1V9SnY1OaYAxGcc210
b0NuCs04UpEcQN83DZaY5sDsoZCnrUy7sDSplzq32rbyxnqjPQdRBx3gfEYPcPgo
mJYv9AB1WrUloIKowHbQGug/jqfkURxliIQbgPifIoJ6jF1xS6RvKeh1IaMT3OiO
/f+VATZgLpVGhYI3h6HF4+0jnoPwGRIZrCRcxdeoos6R/LkZP/JDkmT3qflJHNg7
VnEVWkGXxzEn36re8YaQrkrfG0Z9EWpl14OBhqkZveR3UrZy0Bp6QLA4ivCGPJTu
oSAb8AOlzv+f8GJEYBADx/Lvddx0+299JLgoshwSMJ0+bt/45ZfKSqVoJvbqYQa2
eD7am2ytsvTnhqhO/pjSpjNpVl4nUrxv5UyN+bq6ztjxmwIKE3f67BHIYBE+xeQk
JgNhBWAn/WTmIhxtbD/5WGGYLTNDCiXwR2HG+UQRfJ91PthMKZCw1tDLVYkr5j15
rzfeRolsV6EnQSVjhHg0UmFMRxvDW+RtqTF7IPVjLLeySLyJb4XuDCNTcT0kXhhK
lA5dwNo9UMU28JTCL/v4O0CGqnk1e6NA+9C6zPptzxQI98AmNwi8aRNSWeoGV2q+
b69MliX4B+eNW8Kh3d1VZw5Ax3ncrYFHlGZxPgLO3MDTM6ansBgbmTrPeM+kdXIq
EgAyR7Z6GyN+0uqceziVkZTR8/bAYI7Gi3vQ1kIcd6Va9zwmw9kVy+J8c8QF/ac9
0aucpv4vA1JWdlNEl4cahPgowW2Ud96xr+fak0gMo40Y9oOWNrI6zbcp6KyaJtZw
jLdEGfK5NAhacNg/p+d+UUXuYHnrsr/NrBEiydpsMoF3t6QLVZIpT2BLdQVXejjG
BMwFFVe6WLzJygNsxOB89yw73RnNs1IZ26zqFRbnblYJqGlBdq3/4lr/DZqhwD5+
7dnY680iQfS63/ydHeXL2ZVvDFAD3iWbwFKn2xKjJsVR6mqGqUkUDLqz3mYW7i/f
TPhRx2rAyyA7km6VKf1XUIkpD31nVtC9BmDdGfYzwDrDUE21j+R324/ZPmHWzu53
Y/ZksRDo26CMJzGKOKMyjW/ozgkjebkSB5kg553/u+rOMZEj4s2fcz0C/71TFQL/
dOiqjLXh5ucPaqLCC+i9Kapv5vTQHZn24pwVPuf9tMOdjAX9k9PoAbfxlS/dGVcD
4tmpRgQ/u6EqdjhbImXTB0LoatYOadv2t8avhCbTyczySIC+6DZ3YLMMFG2e/xrm
nVxDu5uT0OKzZUnqYkFTRLzthR/CcQONbGfxSDyFaRHMgVQQAyEicdHnykT/7L7C
dP7cIQaLzoJoFj6WmGqLFnjweDf2fDPB0MXF78zd4viE/iV4W740gqf+hkFTwXIM
6RKPFy+lUPQZ4DPfDX8Vwn1MVZ3R2akkdaFAnQf6sBvWX4fw+myaeWMSBhaEUYE0
TMB8bW4HmNCj/tcrYiYrRlVC/YAL7BA3KyLDOdjfceKppWXBecvGhOWUms++gsAy
6urJu2+KGN2RFdsVgPCPPXUwt+8uxUZ+qIgrUgRs9iXsJAQibknyFY/5Oa2u4soh
9fU9X6847hxpUuQhPowXhfJiRQ/qUdmWY9Cb605tUuai9dFTDBN6FeFfhhGLxAfQ
QDbETrF6tu/NsWl2PIRGsGYCiEXZZLNnOvLM1+CuRqOUQ4F+4Af28abwmbc6+iAf
7fiqV6R41tTlMqXo9p29RkSw8Fv94A3/uAkNsYBy+K/sCTh6gQIh4WnP0TldlDzI
XvjA2gFNKdvs7Dc04Lr7ewAIz2TLO51V/9jc1l0fMMKOHQPeA6gNupkw9rj+6hI/
ODPFmRp5H3HWgAaON0QGg7kJRglGNYy3fkVrBmcxohkn3op2cR7Q8HiM3dcNjAQU
gazUBqMnUVH8zSFlvM6+LNHhTm1UThEaYmGqlBdQUjGQyPCDxrwYlbPB0qRY4yaO
o+OQmsw7N0f86TEX1ahBoEvp03wkHNIsofz8o9y1Q8k=
`protect END_PROTECTED
