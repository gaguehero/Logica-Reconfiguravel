`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h70nG7iSc8Q25X5qY71o1azbVH27GKMViiTJhm0IB5oEE55eQJJNy4o7hkGLTDMn
zp2SBZgiO/Mx/tvEurIkO5Khp3yYGnmL4RkagILWrQKOzDJKfjDa151rSTCPfm+U
86/xgurMv34Y3W7W9Kmg7/laqVh5reooEolki053zT3rEwqLViRziQxhV1JybmlZ
gW3knZpq9YTfg2ZNaM3X0cVa/eompwBx0aUvijbjic1Unz/QgXa2gFQRZfP28JRD
v4bMOH/X4UfQpiAWl30n3VhAckUV/R6z8NVwnKr1vmlmGOoCxykNKX+U5bRBJx/b
lCHktwSxJBhlKUH+gSBxgPkG6olS7Hk/BfKksrbl9etMyw2ZWgeKdpzy0imDd4aR
v0g9vfTWEKCOPiTaCt/H8Ilz1T7V52Etkd4dnrmGIeV2JBm2xIWmQkmjw1I7/lUf
Jl4qduV9txJUP+V6KZnWWVvCHUnFPsPqTGb5enhlTfZqctffPZC+dRcPtLecEOXF
C62JIJx3o0FqhsZwncpSYEhM5z9oBDDkUh505i84XL117uNvJ3hEN6etYCINGAY8
gccitcaYTCXljiHu+3gyrfhTiajVEU5/CvJ2qtXEacmEm8mkWZT6LESTsWu0MCN5
AhvKfubILHQgzc4LsXqg/3pJrpoNJxRsSAWL0LRQxc22nK4uxpxQTvRa76uJTFqx
`protect END_PROTECTED
