`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7T76uo492hs1Guh1dQ/mtIjba28t8opJPdG10lWj/B71x7qoKChBGVoRcYEajEhe
xbT25SlNOu17giORATzdMbc0eqLm1yAanP5t1GVsAf/mVZC5RtgKm1WcuANp6sut
5oTNQMnmkHhhVKUMEG61AVkjAUd9KKJnA3yQwm0MabVU1b5Pny4iDW4AYB1ZwV89
tm4s5I2ukS9bu5u/M4JkLdeKv0IyuKgsC/ytlNx+b+8KcDbZ2tZbvnrma6OjtXc/
l85+NaAkAXaV5otCvvAxETREK3O5gUxdbGHt4Yf+vVdRpkUnYEUpj5yKkz8/eFla
kKv9grHrbVeQ5s2/9v8AO6Ot0LawrL7tl9Ey/IuRwPd+sqPoNpflN1bBKfItpkdX
qBHa4e7AMxdog9jxPInlKdrU8CzuSG5r9aJRGYHNRdwNLX+P+myr2+ZD9QsWVy08
S6xOGvYR8zsg4gkT5SfU+/GRf9lOpNUJDkBaaz8XrJeZ4eLwjSuOexeFEcovcMUv
0dqvp4xSzY2vAcj3qXFRVogjb+eYiF5mo3ebz/kWDXofQ2QALoabmt0kh3K1F/0U
1+6tRjJqdZ6xWxBXZpDtMAIGoqVMMfw5tW7DfVjIK7mLoLc7z14/86Es83R8twtq
TMTWP799Rd929T5k9OZQx+TQLAFYSQ586WptjjCFLMG0ghqGfRzD3L6fvMYk+E1F
A45Qg75zFkcRLioYRGJQDZJkQ/7IIdRQpKu/uvvQLWyu3O5n3aA33mvfkYxJKgRd
BQXLh0EX3OlpuvefR0H8uLgDnt7LvshoCwpvVpFprqONazZhPKL6lK3rEpUNj28y
T4VIY9wDE0XLOVOXWI7MDQt6cnrwA4US3diWXrJjlE+ktzAnESy09S4m5eJzN21U
Pytv0F9kiss1YG3nwQfnV6Mef75zMYUrxOfdo09tcE8jyrMHj5LbGLRmMxwW2wmc
kKWoFhRPyu+poApIAmE7o7iAD8aSF/FoJ7H4TGwm5mONSWGLxP8zOSaC5iTzk9Cm
pESavxBm8hkUDDT6qME1/8iHD7urEKvjcyCRW/txpuaYmrJEdlHWRpao3YRHx8It
un8J3U5PYZqla4XLxEviQRzIelQ1dsLe7j4FznYSXB55W5TslvJhrlh9wquF1KnI
7oXvQqE+ljGPvxqvw9YThZL9Pwc1KTNnyvVBL8KsDjugCNu/fty0eAPS/9CUPOz7
0EXcbpd/H5Fdkgm5p8G7/JinE1OUI8RDIira6RstykknyuMNZDXbvZvqV7cuKCJq
hbllXaYacmnJBC70zDa2baM/PW7b7yIdI691/oAPxUCziDjmPL+qrBbzFnMqHtDf
Wc0fsaovC2kcqi+6YEG10/+r0Pl6KuAa8xldSayw/OIfb3gPxE/UC5i6ICKqGHC3
7ftJIoqzo6qlUaXuIlEDK8RCXgFG8Q1E4XWoGkC2tNSZlXD/XvPOSOLCbdZpbubj
flRZwpFgXfZsdY2X+l5WRoUkiU/oPHPlGAcUn5UwMCJ5d1uIStn8spUD86nHLuTI
i6xo7MYxDl+G3OXLL6gCuvyHqdhqN8G0miBWw0xb4QTcWRlnkGTz1Jgy4MpTc3lc
3AO4lElrNdb03j4x5xNXrHEO8Tvmz0c68nJ7GAhZ+qPGHnnKPqg0UYvesfDzK8ZG
IyhtkD4v/+/afF71KUawXvL8XoOw1uRs3hAPV7qKqVCxjhmtkHwtS7HcIFMis82Q
Hw49tjjY1ImgX+dF4J5iCrzP8BulEqZity0GI3uG2/lrDREbZ59FaJSjG5wnsqV3
91Xn7NaNobYRkoCAjgD60m6QJJi1RzDZkJ4nJAZbcIYW9teNgL24Q3WKFBXukGTG
1MBMZivYZtseDOkLZ2IApexb9vzci+zc4cjQCqgQPb6hiuH0P4X/4aVRjSpGmN2M
mDxZUpSCNTFdc8CzKmZBI4Jm4wvhw5Nu9Vg3qA8IIW/fFIHz5vGCBsLZVwD97HPn
QmFRxn3InzMxCSgIeetTz8KWBo8hUeMv5LGft70hwyieOTzeJRqJ5OWnrM/E9yVd
sw9atchMe+nGeYI1Q+HO9DnZIOiI8J3j6YEfXpb+YJEGXfGHAFcavKFJyRhF57Jf
llKLi6nqtbVsf3Z+2y39OsMfaXE4GBdJ6eMKkRCaeoUE+rjYYosxE4r3Q+4MYHH8
QIat9uWsXzce8AVCm3KuO/Z+TXuzmxWYHGhN3B+zP8l0nRAGDlgpGlBhf2Ey6d4z
3h7s+3ArQY1CeKkjmPeH1KJ9T1X6HJ1ZS/yOMk5RzsuJxcDVWVVkNxD3qbReoWPD
ukUYa1U2qm//tW5KnP1m5sDPkBlUAaKs41faO9ue8loH1OistBNNEB3fPHRS2QJe
1lLmBBHNRwZmYGZEuqR9vVsibT63zlFjxzEVzfHuFAOVbBFwu6hIxP+rXjO8ondY
tjIXebVSzclrvyGaYpWjfSRxlH/NTl4P1WyiuQd+LQRn0efbkgEGnIZNPLcg0X5q
GwkOnglEp0HOZbDMr6fIdrm2REBemUnyuXXSpOR+zBlSUqVhVqRfvfd7o18nz7fZ
E1euwGHw8KplhbDy5y+xbU43Zlyoap9ND6R16cZ8ngDbfItDIzmf2jVfF9B4ardm
sMKzPiwWHrzCdW4eUHhix3eSO6XRZGvp8TUdS4Imr3xvSTfoojsZnwspW1LSg2tV
tC6TnvCAEtkqnucikjrGezERzOhElvrkQFwyix3Teg9Xy0AKs1YVFqDnqPXdC0Pp
2ifdgvCZ99dO+uE/P6EejzLcCNOaK5HDaoSoUHNPUaov1AD9duEKQTFP2KQ2NxfA
rzoMRSqfIdSJrxcT4Ol8UsKmmP1A35pIMn24kcVzDkWa2caaKlIkR8uYKGT3LewN
Dy4x46dXZFPuVzwIpzwyomLcQVdTGOr0z9PwIUPRiidPxfmiZrzgcaAJX2en6O4E
KHFgtQRzmPKbJtZWXbKI83HKc+mRf+cyphz8p4CuFSga5Zt5BrUIyagL0ZFhp3oq
y8kUPO/gDtzScvwtPCxYq3pL4428wg/kmK/XAa75b50WZiOeNyPJKkYWgWhQr5bR
pCXyxF6mfjxdMwTxD6t5Ekzn5XBSOpvdgv3xor3dFKz4QNAL3LKWzZv/NXX6PvhP
p+ilF+HQq6g1LqsyODL3HZDcCK2ZZcgEqV1OYx4EeNnHwaYvwY6H8gdGDjgnoh5D
Hp9OSe3f9CnF6Lr0a3/79jAYuXwW3GfIaOKEIpDoGtgSKcB1qsOoRy0Ceet4PT+5
uoiGi1hh/x+JPKS55SECImcfdt3ufvRLsKLIMK48yTg1U1Gj5qyPvm5x6qfGti45
3HCIjyC0T4q57OxYmKt+7jXzpM6YcdIAd9zVSH6TP1xkLIcRG7c0NZfJw4z1sOkZ
J75UqEd6+LTBqzi83FK/CMRveAeea2u4t7U4VN93TOKM/5zNWrEi0eJHoYVRrb+u
l/WZ4+w+yaM7/126ps//xJF8tsapKImVS1U3bZQ0zJ8Cq+jUEcf5nNy/4GueuRMA
GWw+1BK9i2Rs9eBASLMUnezsxVz6pzlAj9RteGaj5K2MnvB6eujbHH0Ze0FSyhsn
xdiv/GFsQi3ia08x6ubkOrMIPOoZ4mHe5Kc1k724cpBkeRXfj5/ez9PXaj0ILH7d
L9AHpQ0fT9XDyS61/8SdSXcs5X1diSb/ojaCFCGFELNNS4cj+ck9NpHLO2qG7aU5
q+EYk4z+UYEBw7HRUZf26PZplzrPletEwA7hjTyzI9MfvOn8Um4WxGFrqIcbL8YP
XMF4OHkgm2EOQHI3cmuvKgyXJi+FM8yDWq35syReGNjU790OMWUdArijHf28U3l0
zOhcf0TY1MI4N9760EYwUGPKnFX9nBXoZ3w3wgDbvhyywfLR1zh5e2gvo6pBVXbz
obqBSOb91lqDFBCR67NyWOrUHJnWsPEhkAblo0xvczJxygIlNSsrCXs97Cvmgkpx
e45uAIgspqiIfyob8/TUUry0Ho/XkoDPUBvepq8Ohghn+cbLOkYVKW8NNbeN2kGQ
VroKe/pyXKBeUCndVWEogT8RmJUtBVV3eX2+/1ydWK49xHNre39ZxIDCH5FbZP5H
URFi6Hp/ngTuUh74I0LQJr2/rfxDFy1/2lcICXN4tUfd1twWvwMkVPaLpWZA2srr
p0zPazIeNnkvv9Ag1mi/fvrxb8BvCgrfvDsl3KJGJPdUaN+UaBe/gWE6cHnJHIMy
g2t05kCmY1b7bEZKaSCxKlchVCrxSVef1AHsJlRSrlFqf/h8YQljtSCgRc8TJoR6
mjl936CH9hdHI/X7pzyNxa9G2ajX3ZOuRcw2h1OyxB9QfwBUq935b6RWTyN6rh1d
YU+R5JmTwzmNsobgf0MAUj9x/kKjSsnjbzlyEKVh23LwthnbuUMAri94Imz+U1W3
+WNcep6ij9j6L37mazGOOW03vRpWIGmcTZp97WtAEqiEoU4YDk7etgw18sNEbVeZ
7oMyVxZTlpM4MqLrlq1YI8LxhkT8ytWMZXEjMXBbYOT/4kDnfy6oYhYuhsZvaolY
tgVhlYq9SF2Rrtn/7mBf0A0ONOGxxA5p0V4qMidf9XXmt+v7OAEZJUov+fRo3lTs
ivFaS56I74jhNp3fWnZtNljMWJzTX1SlbuBXOPmr8X0H8gEP1dHvcll9KKFnmS0y
s89QjVkHgTH8FwLguxBF2CMk+kDg5HfHtQCYbQSva41/0GG71VNDSZ6F+zT+nHEG
exSjhJjMSdeeI+3NExm3HGE97rPcP7jZNxqzhtrfmWmzM7+bquH7+qoKkvoCOhcy
/KxM6Kr+k4TfbnPK3FW+C6WmpieLuX1LI0YzTPdovYQrlIF8UZF0nXRE+/nSONJK
BcQsWeBGXkI/BtDUgRSnwCuF73ejBAVdW56m7mGqAG48ao0Hkj//tRUwRAsNudvV
cSzsvY9leKgBrgQ8LKeIxEzyH4Hla+pELbXwECwXEFrrsc+mXUgEhyXoYasEy/Z2
Dz7rtmsQxmfBMfq6l1sqH3wbjWyzSonYE11V5eAKIMtMeg5MtTQEZxDHOBR0PgoS
J/WATRCnImocuU8xD+xvzJzKf2LsL7E4OhPIBgbZLeDqCZ9nC8prdXlP82aSoAIF
CVP+sHF/5azb05YWGey29FSQr1nO4ZQVcXnfEY4igrQtYI0GfpP8NnW1hXy/CEPb
Z1eUGo54W8anw2x2lDbbiV5m4b/sSqRsWFK1JWj9VS8fQdNdNHviDqzNSH3MqKup
g1j4cXHUUBD7nHMeS6sqb8QpLiNXmXMi06Om3BmyHv8WCisTe0JDOaQrIu9/qRru
0xFi8C0xuw6VE2v/5qEQ/LLtzrlG78QwQEXkYRUAQi16k1qc/OST1LN7ZgbSCy7y
AjbNXqdvHXDv/b/vGCfke+UJJyKdHpWJ/d9AAVuAe0K1ewCWTAszh0H7uGaSFgFA
zf8yJA3xxoiTnA/GswkU69ijWRU3yAMoKynMmdg/eLFXZh/TLDwexQEa5qdoJN2O
pS6gVOMdwrk69KhGjwVXwwcycGosewnQK+dK3u1vIyAYIoSVIomyR8Wou04nCRcM
npnwEl80NPujtzlTh+HV3L74crhgDw/ney4h/g46XR6BpxGO4oSt+4Y8yCoeP8kI
nwcmCBYieW8VlThzQR3Ri1vO/1YjKuBJvTKRxX4F4RFKf2JzQvjhfXE+46B5Snxb
sGaufbnx/p+dGt9W12buyaND9/vVELt5QQFilClrI0Fyamj6eLYuq6N1ueLWhi7f
Fj9E+EmEBM1XvyC6RnLK+bLnUOuGD4ZKhS4r72QJzmU11MuVHu2HCwFyVEHQxgcp
aZ6T1iTeYz4bbflNbQRa+OzUkREEIDQD477jzPhv28TwzMmeVOVkVyiuEXMFnN46
9Nc1Gi3xJIj/pDWm9Ej6zv2CJnBzLTSOmTKrIkBHGuKb7stRkvARxqoN0LRkG6iX
vEPg6qMwhLlQAHNrH0DBUSD/cQIYhqFd1XsV0iQaoDN8NdAoQ8DXPp5ZXuXj5Nz+
cwwwoQu7saKeBgPIx7bclEHrM4EY9S7mwXViheAPsLlClhhiVn7XzqSFoiMZm17a
oaHEChpxqTqx42RPyMDaihzdKWgiS/6C1RzhS6pxPdeLb7bCzAgtczc1tvKcUNJV
K/3eEaPcYZPOh6JogAQeTBK7667HJhKsDXaJeV2vwXRlarcOUiwOaUdkT3BfUZZ+
CL6YJnFyaEWbsl4AoEpSShSkzh7heWWnq9GB8+tGYzEOPAycYEJuhW/iFHkjTOVT
2haY03sEtZ60sf7Zps8xIRceF6lpAQKc3hNDfeujKFZ50I3tkjRp+uvspmCO+emL
iyDnsmPyTAL7aaGwk/y8Xt6Ps7zGRH+KZlSPvrQjj79IEh3QIN4414g14wkbMG7J
Y+sqz7j6KiyndlVnxoFpH/fNYZvYPKk8xVaxStMRGFl9FSGn+PFHNNuvW2KT2JNp
nuWfsChH+s/mtvJVuFrlU30d2VSgKVWMQrNPDimu+4FKfxJLFA8KJPUGJuXoHyGX
44iuEKLGW7CsBKEPo3rEbbPG5TRB84bD0mu+4yOGJ0BDX6oE9MfToWh7C+59ip1R
72v5/8refaHAB1ZE132HdfNSOouYLzVt9+uNgKuUGcxprNdQM57hAFcK+eOGx8UM
GDZgXkR8ueXWFAVIYMPB/sh8MTpuW8aY2koMT7go/GYH8utcmdUe7FaLdYAB2VZT
JSGg7mijBJ1xOKQtdYkwvT7eQvXYNul1EfFlTaB6xEXUEyYD+8c+InU6mcBoLSR2
/Ru6Ex72YLZcj8qrmXByG8wgZG8wXVjzSveLo7oFvvFbpUakL6PLTFH4344lQIXv
WEN4NDsbIaopw335gtuDOiGSDgzan003LT1Ay9K9myrMMCDB+9J3aGSeT1ZX4Kjc
xofGgY/Q7PFFCOX9KPtW3+NXAcgnEjknKPNfF2AsmLneAJepWVmKSMS6c7VPYcrD
f/MXHcAMFtjb7QpxbxkLEdWwaccjg8ezXVsM5RUDqdMVBg5SgCmWjR0X4tfUtNsx
2Jf72SIOpWNiKXJ35eZeXLHjR4WSHZnAMpsiUxmlnWvUQRbqybkytudPmDt45pch
kJyLljGl5A+xWgb5TzftQ4iC4YAu8O3alByIfJzNjMdCwkj8b9jNtNRx5/PPs0K5
SgnexZ4pCfqZga2JUZb6WNpfA3Fka8FQK5pNbj2G/LXqzof3E8NzXG0+IiOJINQv
ZsQnUpfV5p+m80aARYAf7EiTcTFkWyrPXgk4Jat5dY++sZEeRqX4FcA7het8ZT2B
Ly0WJ5on1wggAd1f0USY5gCXCvYSmYvvPVfgoR6O3pnp65PwA+vDD2AFPrgjgcyY
eVrs/vXm1Zge3yQCDyLo7Ba0utjNCIj824pEtCy+d3uay08vOZFTyVFxEdewzXp8
ebpVZXTDknq95gJLiQ+iQXuEsfd1zJMdzDVa7rb6SO8HCNqWA2JizmhUuzErdC5i
+okLBH6egDVx6LEPBAulmNRJE7KJcP/vpWbqbjYB98FlNdQPzlCNe2S3525FN/2y
8N+sUELxXsY8ssvzKIXSg4T9pvFlti2wokYWN3bi+1GP09uDXCW136/XDVanxAkx
EeqNjDBEzmrmlMvUHoZeT1mKx1dP+TvEcvBx8C0vB36qc/UPY8naAPecCvKuIA42
PYk7kYZ/A5Oz2lmdPx13HVxsY/TFuwHRvMUJJYfcZ+X7FyiNp1QZ9Ws+muoitghP
ioKdY6wnG2Npm/MzitIKMTPRQUlzUuJjYVrHEOkBKt7umJvpvppTcbz+UnYuALt4
3b5HNhoT5INI7oKGOSMwCxzEI0MZYdE37ucE2BYIR3sd8ofQ36r7QS43Lv+gQ8wA
MwsoV8TXXXLpQU2FtgKlLIZ2kLMGkchw5arVnLKbkEzsGfXqSDnR1rsmt35upTl7
276gkLIxEoU7jBZfHKC2PEJ6wdsxHQk3aEsHzFAv+IGv3kxuM9AtAeZNw51GveSM
sTfYMXYSOKVJ/5NRYFJYgxzWkBY5+BMia7fojviMTlFO1Y83qwrHfgGojHFTfl1r
UAc8Z9Qzr5HoBuevH6QPxap2tCozNVeNidBVhSq2S8VSoV9A3VmDvT8EEm8xj6Ch
MqirEW4t3Pu5EDJbA4JVwJFiZuXI9qqy9x7GHAsVYbY+ySz4iqH30Z6gR0GM4r8T
S4c1rjHEDf+Jnmo+0VXKYf76/MTPb8F4OhVgyZUe++sKGkEE3DuZruHghAO588Nd
5Ar7sIBtJLVSGt4JZzxAHS79GlWBKtUvdkVXrhpToo/Mz9OyiKHMIxqLSb3hVeD2
RjO1MlEuU7OTJ06goLakIZDLKcbzGGwdmcsyGQMGodurRxHsFyneqM37f0RnoWOL
wNOi1JmnejkVKoErqWitqU4DMN/2WsVm2j6ien/kz0wN+l0bA+6pqbnawmYqGhuM
Gfj3uNRcfIssy4BAyFP1bQWPd4g9ciHxc6Wg85kssBIW08pE2gaPA3FZXJFhD1+x
OBPzvsFV7e5542xGV7TzcY84Moxi4ASRLqXfESXn+Go6mM4qa02s6G07VgQ87ZDR
js5rNJiDo7qcpD959JbtIteuNXPh3G1rDecURskrdzGhpXyykg/Wg6z6tTEHTznc
sZzixaDWzJNgjiHotJvv3yRQhQ+TpOxEaywEKt+GXMMuQE6zBeuF4VPO3JP87+mX
oJqAzyoUz+mb5uGxPQU/QyPover6tG4fCTFuiO8kdHGeV8AfdexZoZUkIN1UlH9+
MY+MBVJ/b+54MwOtugk7ebtlvrLC9S1irQbd5OEP+FuUpqXjMNGf0l76sx6ThyIU
W8LxRXB8j4lC3TeCavp15pSE8UMSm6st20E8v3gteLpM29jMNqwa8+oCZMWfuUWN
TbHX3yRcbEAAAGqZVZQGyQgRo/fKRSDYsc1NiMceCJAAoMCS+xxRzwmSbB++Mo+9
6joEa4bGv4QHx3KM3mqIuEVR7e6ocjkZCOpXnaT+6Xlt1wpRLCMOHM4TE2ylCUSe
FGlZrJrco7Z0DeJ7JYF/Ak9vUhxFZ86apOXaW4qBVy300Cjq6+pzMH/H8DGotEkO
XEaim7oj105cMVqcEOElIRJJgbN1vlAi2w/FX2T1gD4rFIrnELTUfrfCcG844+yM
o0eFjhEZcR1Qj0lVPAyy9J31qH358WeepLCUnSDecmriUJBRowYvPrPTMD+zYilS
DyBrijLDfAhtXFo3qLWzP3QHXK2PXNz51sYcpggqSuZXR2F0HQrG981EgjrJNRQ0
NkDqvcBfQ3qo1BrlXrjFHrlSRtlXJCRsv9UA24TyupA6CHH3o39zco5/Ec8TmsGA
VDWhzFxYhN5TPmpZ0gz1Fpl0rhwjJw3MFq7eUxrwlD2WsFneHHN1AkKJ3ji/yIwa
ZQR1SyIjHIvQHbvReqWkO6+vSM+i9hHrPaGgKKwp2C0sykbEum1LbfqFmevUZTZQ
h5GTDNQfqVhmMoKDoI04xb38QAakOVnfFepKwygW/W6n30cX2aQTywoWFJgW5PYX
Bbn4CKkoObyahPNOTDUYeNwLBe5AVqViLmgKW8AnctBx7fyTn1OoffvSviw693hO
7MjjvC79a+Wu1TranOC3SWC1RNYDF8e5BBx81FJSOLoO2/uNGHpb/P2xwBeuclr1
V8qbJmcMv18m0dIp/3rBSgBfBcDZLk0iL/be6F2TYjdt9KOzE0xjsoP5WrhCn9hE
JKLjokMaRzSfvw1uTsMVhHsv8yz3P9Q679NUqCXCZDdJcAu4LVI8Kf7v1Ox+IfvY
ZQ3kwCWVyPn/qrW0Ho+6ron5ALNCWjvzY+OdK+cF7vkb5Mz/Zj35sOM5kF/nSno5
ugwaXEqL8iyzi0liEKVJVMRh17dnQkM0tHCNqkHZqS14k5MFGUrv+3KOrU3MMxy4
TSNtydm/hojf5F8cS98Qv7tRZ2KatOlh9NMri9x/q62bKpadoxojmjl+c5qp0opl
x6yCz7we3EqsdC5aLAtw/kMTnB8ctilWhVqXFTv+o+yMU3HuKqgDsjbjZ2heh/7n
fNS8BpumbwrqYnacSArXv4I+lf7Ast2WWUP9V/0/VWiSmTQ1szv8+5AdqdgEmWKj
DEugEZaSTbt9v+/saNukFewwR+SE6a2R+ksbE3+aq7QXx3jsc6tjfAjN+fuMFr/q
iKlVH6TEyp7iRpWQ5d2RjCgLFbiPGgkCptnQ+3Vyqpz01/833tT0I6LypyhgfRdF
aUYVUS7nHZZN/Emq3HnxdurmI5t+TalYTvCeflAs496pR/PYSCpy8Nz/TwXZVRih
gHALzv1dX5tSVDiMk4mPvh/uJOdyrCnBWn43prtrn7Dr5tvstvimMGGdy/eDXgQE
L6u3gHQaTjwG6QUNtz9MMTq6NU1VGr2LKLwlG2gXzEhpdxWrPQoww+RTmzCHFUJl
3853TLtdUkZzUv7eHgYetkDQgHFvDIGSPEUDZkT52Dg=
`protect END_PROTECTED
