`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xDzJ6eo4cU4Ls+rxWxGPfoCqVJYQrfUbu2yGjvxXUefnSizAQLmSEF9+C6A2ggK
nqpA6xZuoGaU/YPv62PhFyDBDpmvU0XLF6RZQWxgg1TkaR3MpUy92HwdQkiMopqR
s6k+Qx4Mrw412wUcwuOEOc4Z9Dih1MCY1Ymk60cOry8FjPN6Pn1/S8YBVV8GQOF6
q8Ot6JHyrqnMN7Rj76vyYXsTG3m7wIM3NJd9S6A4f6u5KkxewxDVbxGlSeRP35he
VhHLIfJOnXk7y5NOCyNugZrzKIG048jLB2+QfwPKXWpfT1htKCVvqF8qRxGGFqMp
ocWDmK9wKVn4MJUPPhuG2r1rY5WEZgWOBJQVyZWgewkk5fioURteE3eC+LB6qBTD
obPgGcW40CfXOQ1xvezDgzEv4jJfm12v6WjL72U13K9cV+niSt3/B8JLq+wu0nxp
0pQ6vbIdJDgxMF2lB0kSbcm4QRYPp7mnz3e69BjRpAe41TedloPqj0Ihz73PATQO
T+BvdZORP4J7mIIr7NVSjtzmimXXT/Hgc+M4Av986SXsoJ1y2xrBEhIRFHY1HYV1
6Xiq6zBsfk6YTBlPxsn46ajlZS3ALgu0fp8tUJNZtliHz10/d5Je8mfDVOZYo/C4
5/bN98uXdKN9qZvLqDQSpuQHATIUu+n0yIuSfIT08CGZNqyjoFZJ97q6vbh/Ai/h
8TuBbMEIPpqYGRNcnTLuU+y5Wbu2Q1WQh25+UWSualAQLwpUWuUBEjS8ThiNHPvB
PNQ/JD5tjqtoKOa+w5eON+4F/fSfR9nWc8hSbRtBxAPkSMJ1Nipe0hRbFCLIEwmC
IQFa51x4bXcCdwlSIo73aRTzSueg2a7EomDoWn0byqSRZsdp5wWsoCeFzH619f6q
NJSs7ODOSW1nVzamXCwkfgYH1NfVZO/NZM9neuk8GmxzW10wyUGJJBeGEIvQd1XC
x5bRWi8iJJpKF0N2Tnqmgapqx75s2eST54+GofwMtOHbxt+Kw2WKY/WHeneYVSsd
Zky4s3/v1kTR9zA4rKj/o4h/xHh/T4uHQOzCj2CYnPrm+mKnUMKXA/6L5BEf3SS3
Rq+tnyGtu06dMv9LTpUbxCpPneF5tTsVDlCmFepgV0KLZEElQwtR2okpjUmFe5PQ
nr4DfDW1vK1iokoN4HHysr2uZWu/wu4Mm6SU36AgteL6yryrDHvHyYsrAKXHONnS
0CJcC1/ovtQXmIWW/nBllHILz1gsL55PMaaaVeipTkhB6NPjRVw0muHeNdz9kEe6
yVQORGW9zm5TNu7E3v9W1ESXOHMDCqF0TGbfunvKei2EX4ISPek+nvwk16VrZXml
y+l+fIjAHMgAvt1AU8Ew+FEbaB8upTUupa5qPt3zLwH0x+ILkul7ix/E2t3hx607
QWfV39Q4zJSSxakGbMOEakIukJKpQhKFhL/lES2l/XZVoTEwcHcPt5bnhTEyrUUT
7Xj+DtwykHxasjDoAfjAibz0pnWnv8BO7vb6foiNamkARwPtGsibe5yyRQzVLr4g
yndhnuLoO94jRPuLQLoGKjVxunV5EJhWEHehk2PFfjffVbnm3K6s8mve0kJTWuwX
DmVL9/hN88GbuuDBq46iULR3+6VJApcE7zp4d4F7zxPUZnSVkEB2PSqhYJTQ+Jm6
Cl8hrsxs6RYyPnFjVapO9XcqD+bxBNit09gvJt5I9ZXG8VWDML7jjaVb97mCK9iJ
sBX6cqAjq8FepiD/Rn0hctdwkxezqoCWI9FteYkDYy0MHFwRMXOzKGMOopirEFkz
7mSUB2Dlruy+R5NsCLK9uXObh36ehYE5ZqU/fYykaFRqGwueipa8Tlo+eJKEM//v
HB5KNI4ePaeaSdTwg3fshhtkQryqIUC65We8UPJYp1P5DKTTKPpPJyVTbzaeoh0Y
EZw+5NeC15owQp35IPG0Q/Uw+W4COPB0enOHtnwizPMYNpYZrM1mKnv1curTpUBU
4ugGw8n0bC5Hf0a06ZaDZrBLxfb3qffLBeJLlnUoZt6mVf5wr0kUGiqIPPcSS6u0
aqDR04wTarsYgL5h6OLMv9eUthFUX/Cl4wauthdFIBe8qy04vhUXcb01WTBk6M+r
wIY+N5P7shspz3vFMu+arMLuktVCskXT/O5lnpRJ3FC1tzM+xj+y7g/C8+q5aS94
esx2q2iMqYIjBhcGi3vT/tz8/Fu4aQ6/peNtNyNb7Ca6nRTa+f/y4ZK/SiXiyRs6
KjUn49dJkWeKCHopZ7mWRwApaBSujCAkrlvI+DfN+xKERT3kH1Kew1LgGBzHrYJY
hbKSvQwfnqV/BnNXaXC8A5BSsjPL2Wma8tFzSEOBdFcZ76UykuCxVgRdLo5i5kDa
BFKyPjADr2FCuI+uTXFTJolpHSkcVKJaAlSpNSpeWULe+veL+SgLpJe/Ejd9fPub
6/ECPcCYn9ZKjP4Pxcd8T2gTuZKM/yIJrU8pjJzGpjcGAm5aOO6VWverDkYlq4a8
tFEocXAlCZS9FbiEYTJBMbH4W2aXzMjdgcAKD94RdeLz7v2cs0nPi1Y9SbFBbSp0
GOJcNhW0uxqWZTXMkqvDNWQrk+GNUq7+rh2AufCI+ZfoBxTZALuowyuW9NiYVrVF
r3njbEzQZ5KxrEQ2I8h5Q10+OMPBYurvI7+5ZFbDtpByORlE1do2AQqZjzlfMCOJ
q4r3pVmWnd12zy+fGf6ywOzn1aCuRJdTl5KZ24TsTwzP6OF00TKYWrBpgHaZll5v
FOFwOByFPtiyuZxdUBNT0VrveBkcrUDY3YTRvCJ3HdxXHJGnCDjKPxkjl+G0UORs
KgLB57aWqLak+JrqksOw2k8DNbzsH41Pd4JzapxA/ai8hh3O0EArKSNdrYl/0S7h
7Scj2uoOLdTyzGaZ0fpC2vgNbIceRhKeSZUZ/3nRovw3aCa+9DNTRNifnOXYjHR3
Pm1a8s3n6m18mFDbC3wXz2tbMqzgEYjOSy/Ie5dhaXsmY3uq0GRZzN9tfZkqmDRj
1ScKhB2wpf7O8x8IQqm1bHJIVjf1odqHWsNTvyQlr4w22ElplIN5w4VjwNM3mCUP
uUe3vJgTtaldjecFvcf00tQLwCZIMo8fgXNOAgAhDIE0xdK4TEmtLcmUzrICW9ui
n4P+mXOQbA0BLwp/4pM+g8OCnaMaG4NDTEAklV13cA4KDoQXjTqE6P1tYHJJbPfs
Nsm6eeRSNsnZtuLGjDeXNIikyomd5gWOtJl2GBDAUnKHeXFelURdZSRZ3vLBIgit
hfKulACgqboI5libhQGlXWyQnA7CJzVqV30KZRpeGlM4Fc1YWCe0REik0jCApfsS
mejaiuBlceCXKz4rPcX76k7NLs/SqRrgRCH8KRV3dgOiQvGHBWVxBDuN7r0yk9bl
hy3FOI/P2Pol4nV46tOmhLX+ztc53XkomqhTJrWg+cJaugPlCGlrWqMrjoYWbPTk
A1+RQVL+SRZzFHDBZ3nrwRsCmHO8PkPb4PyKtELWwd8wq2brlL+jbiAtfeoR4YBg
wwDnf2jEdlXDxbRxHaqh4SlrylrHFVFkLU5sTryKM//fRPv4mo/w++4vmDpE119M
+Y9btq+Z5GglAp1yUnIuKhYcRFss1e1ZRjcrAgNihqntm93cLqOoFvn0yeQ0I89U
XL54cfXPl+6/gmDM6WbRxFHWGUEeZQigR3N6BaHPw9BeEIFpZ3bTiDtAUsMg6vAZ
/ngetBQs0/wX6rbN+ZrcmR0/ng168CPM/HSkwRqrd97FTxXA4a+LwD19W8YEy6/b
vxQnK0CPqTwxL/lIL7zt5tcaK7FHrWtUwqYkUT6ecq5nx23RtaYlwcZbhbJ++irm
4L4PIjgoo2C7Szq7albZadbSpQJOE85125agef5vni7oTKLpeVinXstUlfZ5lHSk
ytTu/c0APGAo5B2/yl7CMsGBGmx7tZvSZLGHekyNVptKlhu+NpReRIsSOXlE23DQ
kHm/R95e5j/YGxaKgS37WmKwzBc1nHGUxCVTQrB8dPJ9P0ZC1kr/E8BjoFz9m+Nf
B6ZEptPEsVX7FnkmRE+a94Be9w4ZoXNEqMo64Ix53Roah04LrHDOsTkjV80NB4Sb
GZaj1heQ+KD4dXEs/3YkcBBm3GAz0yo8tdFs2RMyJTDPJ8bvNBltbb+y9rj9adDM
IUOdmCm66JUSxujNT0PeCwunwMGuM7TFymuyBJFFYoVexPge2bz0TgU8N1d6HouR
+ZtliskFEqBuJPYZYcTDeaMMX59HQOGrEC7YrDaB87YDoLB6YQEUqJ5CItfwrFhs
1QvMX/AWMtLcjBDvIbSFo3jH3cosR7M4a5ZJBrVr/rWe77airps/W+bfkTtSDM6g
Z23igs+PoYKOXwQD7wzTFJjNNGeQ10+YcBaZXgzYvyaJNW33cNIjWCDwPWqzQH+L
0+X3mKjnLR7Fi48cx7n239Asj2pU4WDb3LGCoUFvCfCn3PlGyTUB1h0G6n6BmrvE
VxpSQV8fppfrm0X+Gb5dPHZk6+kZQtj3mCZDTEMYXW5yKQn60C3e+YVQUMI4GwpU
q40fOxpjH7IE0AuQDeaJa9fN7CQi29ywKo5fwabPnIUK83gyjDu3ZsAMzWtKY4wd
/2AKTdx2RusjhhlyD5m42O5Ub9bOrxrT50HHOj9v0kMJ+JqlIDQXy3hR4MINu2jg
kM5gYzzXrZi62gdYJR3OjQcaSleWixaHhkrAIeYFaP+iaG+1jnNIviacIliQ0F37
AmkiNZjWGeBdz51oyo4BrntHh4A/QGEol0/aKgwtQz571RUN7BHWvbHPwO8JQ6B4
0qN4XxtO/W4aJQW1LR4E6q4MsDosKwJY6zrdcNz9nNeznkou3MvnwAt4+WC+wBaA
6glAQZtLjq90xb8XzQdWLRhN2q+eX0EXjdk0/XvC3dqXE3aheaz08GcTjPIx5Z4D
iguDv5YNVAvqGuwchCaSZ7VUZo4U/3ntA40iY27Cr28kW4bAT8UjQBZa3Fvb4Feo
0+/rjuwdRM2Gzrn8b0Vpk4cg6tjXpdtwrR1bme+8OFBgVAGpGZt6e6UgL2wzrYjQ
CCq117fPcyLGGba9k64RKtPEv44OXr4kf0Ygyqcz24DxX4spRcDfymerZ4Gz1/id
5EddCoRj60+y6Yuk3QFMClkoafEqsuoJWC2bkuUYtAypC9kcGjc6K9qwPF3A3SP6
F/o8+TErKK3oKVjk1rlyxcVwyd/EexWSTUJrGc7vYRfHHyaZyqvKoP7amMeRQbUu
+klhZliBFkHX5ZZHIu45UzUXBNw7LJ1t/ya2CISVs5GEh5FSrPB/fG70xNdBiaRg
776iYge+eQ7xw9sciPa+n6N47R8nrpBloPkhLWxS1qgLmbZJWV8bb+NSW1l3TZw4
KpyN/COwfjHRKleXai4PT34zMUoPXZ02zsGQhOaFW5yiTie6xNK3ZUQSY5cjimm1
kVLSW6hY4FfsaldfMLQ6oxb6lnkiG7wSFJAEfaZ5qpQDhjyrgBlIret+/ep8VFgL
uzPc7L4TR+P6uQw7V06NNFY7YsYMmsaisYsoyix5kI8asteAl/fVfzNTSCdAy0zM
MJgRGek9g4StYpKTz/eMbN1uHr5T88XaTVVkyP1FDLdYY5i7MXhiT8CGa1s1drdh
rA7phrJI1lg31gIU0Jofs2WD7t80RHkwIBvycHj4kZwbozGNspV3bsKHuijnsxxS
gK9ioC5hYKMTAJ/HljR+M/CxSPwxZsFDj2YjAIj2rdM8f/4mQrjcmHz+uXEWoKpq
nm6Cn+m/JNIEmoOdgaIr3MdNPXCMgqzqd1fVx4eudnurbxKM7/BrmGVbZye9gkM7
rSk/S7vaDhEsMZc4HRMUbrHpaswo5qWT33VQTiwz3mcxPvVwEzTLXv+SkGqdCiIu
3F11DVHdecLFpyjy57iVNGod9sXNHLk94ypKoOowM+UmjpptHn/es3E5bqSm2H6i
K+gcdlIpaqE8KRRWdW60Dmnrrm+hc1zphg3XTOD9K7vhUTEdCxl9+wf6wBM7lFla
rLSoesSWd/Jk9inQsRYdOoHi2Hv0wmDcQ/M+V+8AJoQz0gMGP1SARKFI8gzb4fgD
6lCO3euyu8T9amnNHQlKYwGESyIM2X0QHDnViQ/qQ/dtG6/9ic27VglKo3ZAM7e8
uwvG0hrw1hGCf71DdLActtEA9zoQ+OIaQOiYjrwM61lDimHbFqFyihcOYFrNxrIE
i4uiNEz7W7p1SY5NnmwmwTGXuX7Lmc9HqkJqd8Li8PBt6ERGon5etaXM+ILdzyeD
+6UaR3pKUzKdXHHXd1zrnW1QcH6cn0uR5DIqVOZ/7DkYTdYW/PV190C1GVeKJKyR
UeJV69vdzdVYI0/xvBCJHRiuI0SWvE0FQ1IusbUEeTaCnhOzG2MBTS9D0jHaL/Ry
XASDbUCnaDETkhWFIbx6X8RhnMPviyOiVxJ48vDsrnq4Bgr6Og0fMqd9TV5f/r/C
enpHp/psVaMm+t/W3n+dxBm4EJoRM8t0b4WCyQizbovKX3uxSGyexZeCoUag1PNs
v26n3fGpMujxI9yTosENhdK7viuvJqS0+ibdYnu79xhBs9YbEV6/6uiZAW6aCNwi
jBOokkQx88EsqpJDgQsXMkay/LK2Q1SmMcdWE+W/6a+PSnC0VeCbI7BuYCbW+LkI
9b7nb31ajBaURYMDnbb9uRl/dBTFh4CSFNBismfmyiNExWZ6fIhXDWeZ+gzcNQ+r
KtDY+4/tZhYfHfdgzexOPbHjXM/la6pCE5ilOTGZ/n6yTJ7QBEyzt3R+uvuv92vF
IJMI45jfuudEFv/JO2jN2nfv75Ertvk2EwaoDnXaehomdqY6WbA3/drgii22caiG
NKj/5KOa5OzdJIQddj2zVnTlqYjbMBDaeElc5uSsGrA4B1BVqiFwnN/4hS2gODmH
D8imymtTZm6kCVQR+wKDO1gtA3fojPvWfGWLaNsXZh9HAqhb+ieiHRX/ubpWnsqM
rNdbol8TCMWZEHeuzt8MAJ+KKuT9lYjHvMiL/yxB8ulHVpOwRAG9b7qgmL7sPtF/
bPWJ1G2mYmASn2/an3iyqC+Q1SB/HVcqWxUc0UJklDu81CKnvQa0ZiuyCiq1AABk
73KRXv0XM2dwCQbdPwXN3QuIQF4EiSu+GE/+9dNyz0hxp+ubmxCxAusvMVvnoE3+
1jzPbP7lueliiVhGz7QGepAf7FRyRY3tMjo8iTjvfq61FuH0h7nVkQH/B0jSLr7I
BlcnTw0cb1kHnQJynNkgjPATrpTgL/k0bB87MVenLH53KBTJ209+/vb7r8QHqdr8
Yptfm2xarV1qIvhDB3vkOf25mXj7zOTVHhMkzcoxlwimYyDSO6zaMP5jBu0LOstE
zngpMzdDm9y4G0Xd26Kbf7iwazgTLko17Kdmljy1YBCk2AhjIqz9DLjMecqgKFka
Mxc+YZ2vHg/SQRZYs4vEoRxzOs2RsriyOXSxq9kKZOtFdfGL9Cp+jY2Kohf6dQs7
obFLnF0JF+CVbOLzfD0Zw8jA3AjgxfuI1XS7/TLs0FMM9BO9bOSqFxI2u6/zZkS4
8nRpyE+jnRdY/zr4mKbY7L5VZGPhI3+pmUy7oS38yTjG0OYZJx9pNeJYjlr6y3po
VqmVPLJSkZO8tQTLiJOeHPh3efV0yruJAgfOXCD3c4SwW90HWxmZ9OdVP8uQFjyd
WtVMr9HbQCu8QOH41or3/Jxuwzioj8b/gMkZY4M34etS2UtcwMzP6Gv4knlWr7q2
a1UP01yezgk8FiB/NEK4P+mU8rCSpcX/bvD1pnJfCKnzYFayFwHAmtwH8jR+Hbie
PSh6MMqShfcBptlhDE0i387Gq5eiFPNdM4XFe5dGzxjhxy5FMtW1mHsWa3S+p7l2
Hpgpx8NrkDeJbOvpJOLDi2N0WCghxO0frsr/NwfNNEYTVTaoYQsJ/z6L7hkpGOR9
3vLIVBK/RQ22TmANVBRpnMZX1FmvK4hdqsHSpxIA+7eHxRk5PwhqwVrF3c0ktaKt
NCGjziKqp2dZroP6aqOuG/3jps1OUU53DWbB7KZVieM1tYE4LXC0hk3w08E2E9wn
/XxagSx3o4sLLWzZ6aIgA+oQnY+bbDfAbmIZs3naIfifAabQy0FZV7WyzXmPd32B
4A9ROXelHfuZ+IemAfnzXN254iL4nkLmt3RdCNeoMiE/IBii0e62nuyJXz6UtpPT
5CsVganz/ncAQDKoBk4RZlzOj/rr2pCTUMWXuXmPTgvE0YppnSBKEU3rhAaoBL0f
fR9Nj6PiP8zbFKxnK/+c6MP3yLbSXNyLcZC7CxAzG6hZR85CC89HNT/6XTDjEm/n
mvup4I1qmtpypgCnoaul/uSpDQvqzrz49fznEW+Fy41ORJodTtOkRJYva7Vyzm5S
K0v7LfJuaxToflH5J5YQFIx2qfhAvgY54AzOAcKAxKlwlp74vS+4hSQRyPh1R8DU
fCh1b/o9tPBYi0n7bRahPzq2QIdE3nuHO0W8JSWFanQxe+zlRHQxy9rh515zvHtA
bQS3hQlY9jT8YvP3LwlaILrGufJkfu6r2mdRZGqEb7KwVy2LIoD7J3lOAC62SEky
41R+2hTBwATM+V/aIph2tHpWS2Bjlsq9Lfw6TQCUvMQ21H5G6+atcqJUHtz43QA9
2jRrvxcSrnkjo4nFdRNDbWvOiWNqrQ22gyI82p1jIU6rLlTjnxEdMTD91mqS9E9W
vJDh75x9vx1hfXEhNdD3NC/vrI/Qn3wXZqeHKAy1KS8yrlxw8m6jNunYTTHbEYHc
ERoxgt7lW0oKLbsimJ1a3Bu3ywy/BlWSHY2b+g6o3LjhKG9xwpnz7SJ1w2rBrQn+
in0ouKHRzNkbP0VQ2ruaknnm0AZH2+ektT7SCbazbgXDMpPyk5MSfWX1+YLaMnkm
m+69axGfc/vmsCiVJ7i0iy1lxr8ejkZCqtD9tDQvHN0=
`protect END_PROTECTED
