`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ud57mhvWmkeJo/9LCdTrmQd2nYYiTjgY9gAxGS2KlHcBvCEbxaztxW9L1gdQVseC
hBWslmrFSwYlVRxQt+8qRF6sZlecCUoDjqf+a/04KzUKRu8wOyDT7s1DzHgkPZB5
X9HB8LMhzB4Y+DktDKkDnKg8fbzAs9Z+K7iVID6Ssg0DO8Rvfekqdcl8Up2aV+61
8kcwZbM4dHXO78bpXQ8si2Tr/ecyqFEuMd7NshWyyaeApYCclAy/V4jjFLQrpwlC
gG5doBPWBXba/SrKofjBZ+iY/fYxZXfU8/l74c4cNTrARDACzvnjZTx/57L9klgY
ula6LKZifxthBlogTEGLeDmDxFOuy+kItnYiT5psobgPKD7cydTgjQ2kOAYNk76X
mddsvxVJza7IJePMdiQD0fE4dH0Fc+uSjpoyCY0Ubgs+DEI2+OwzAcG5fGKzIDwH
UW/mT4d6WQ+dSy2dTFpwD/uii6ACrUA3P9id+RWrGbXN0Rw4yf2N0YwVdsmPpQ2K
+Dc0qwp+q8kc0WJmATBpG5Pmt+hEVNe4izWrFtyWbLsvqZkg/lyIVGGekRt4GXyx
F+8j3ZUYOwyfw1a01UvNsObqzloVsrmRM87FBoihZO3v6fplfK0LkgGZuteRkpjZ
zIV/gd1/DIveLB/+sOQKqCNvmqEBI0Abqf6NnSnOgmyTH9HhXzdmrDli+yFcbK2c
eezifwRsMTL6jNsBNDbrlgnM0/4eGWM8FWLeKVFyJ4PK53emqifOIhjHuhOQYw0c
m54dD89Dzo/R1qcaTXFE3/TaGFc7qqi01GxuMaeKfvEWY0G56nJ7c1dHwnDMVoGQ
A+VctAmFHk6GpGuJfaw1D0XmfNmlqfTXBB+9klE/L5KtCOzXJwB18p/QNi6VTC8c
+Tht1hdRLTgmivfehh6MBYl6Q1kZRup1GV0no15tuUTHtudx7f48DAb26WHWWfBm
fBWogngOwk4q07RMN8WWfi/tVsUZFOnuBfYs9VQuKEGmtTe/TsfDVRE6em30EHRM
4gv/179o6N2Oc9ZYwINCMN0489Bt2t/yUZsqJL/56jJbTo2QlfDB9xKcSRnHAPm9
axzWV+z76xN/EPQfVp+f0fOHE8BoX3ejruXSkcbi+gop3/CiKrQtJI4TQRGoSSnb
9d4dOoyWt/398YwbAVT8zIMkOIBJsKno2HaUDZVrI/bYmp9h9BKl7TJHEgmQpH5/
g8qJ1s5m2/k2+LN8tUUm+s+9qLrZ3NJMRTBLHaLaRxJy2THKwiYnQJSK2gEyW/5H
Qv99O/4n7FzBBFbyIZch56lwRfcihZ6srhmUBjduFySbqfpPHokHwD+ps4w3okoF
ik/FFTYT9FDNZkA/XvMUStIJhkFsQ6zlVzxwv+a7usPEeKQEICqHxA4vMxRnzM0r
lU/mrUj/ghdPXntjzkBfu9Qv3+mc1kG6m0vfIN9yh//B3R+6dg0HXbRC7oOm21OA
W23lk2CR6qjIGbnm3qVpcMECnar/q9Gdo2fAuX+iqL5/PxGOb1ScIC6wglmq/7jx
NJbjdm8nZlvjLiAAu1PMXVX6db8qabmDy8C6c523kVmJ/nm+d4ZVruDVahFo/EA5
n07Aqi27LlTMwqNwy/SLgJY6W67Te3fWvK//wCTnNJ/RYjwXjslXpgd7brxV/X/t
lhOqPFzyFK+NDA9ylyf+LQ5mbdaS2K28tVQ+stuPLkNZVdpQOGw7WxZREHFghO4+
4zP+wuKy93hKyqpQQKFbVga+BhNEvVW6xbj9ysZR09RJ5k3+L42FJhqp3UNd6C1a
BSS7XQNR/8kUBwMK2n+6zCpW4TvBnFLdUaxJnRfDUDxVbx0/2VxvnpnS7sl36Yf4
VMAtzsXsLyLYHF1sXW+dpd+qncwv+PjKpmtDzsnp7fPYRyQqrPPmMcbKNcJa+ccq
dvUd97BEhpOAUbFfAVt4ykc4Q8HEFG2Q7gw5naBv1+C6wTVQFFVa9KuYryYgElx2
iFehjdkryA9Rp/W2Ke6pKJli6viS2YTy1FISxq5vlW2QNohV/UsgKvbPn8XsVqoi
lCm9YbZEKHP3TonMYeOuoQ==
`protect END_PROTECTED
