`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKsI27XO5FqEAm9WiOEBmUbEWhTLY361d0NrBPItAcGVgJttHn7sEwUuB6r4qZG7
FXAEuP5/XFY1qXbBjJltT1TyKFm407riFD2kbK6xQXlcXakMNTast5xK9e9eHYVa
ve0Olc9JxqVhe1Qkyu79i9Khfks6NsbDDaPEnVZctXgd5CjfZs3tEKv7KctkGMMt
xADHr8E5V5zq+eTOWqIs96NgMg2gNz8yFwV1ByA8fyUi5CJK3e0NDEYj7KO5Tx97
MVwcFJnYf4kpqlJp/RcF6r06ZXWT09Rz6V3T0Pxys8adU1YYfC9Bfa9U2JKC1HNk
5hzh4DUvyb6bCB3m9h/mWbloEyoGOJQ4xirii3epPV5/JzbCnXoBkS91u9/Ud8Ik
XhTGFMEy5Z4gdgIqV15QcDBuYTQkB2dlBAJtHPOFDDtCALFpJe75hz7EzxzsCSYu
d2NJQ5zEmiSBgfAwTBjkSCgJ5p6jD6rpJxcw/GAE/qWB7od6REFT8VkueC4Gtqg0
GJUAzqvImpk9P/G73pGg5Fh6aZUWvm8UaVlvHMEW/KwjKTOGuk11zKMxkSR9ibGR
CvAhZXSJSnZ6fLkvmhC8fjvcb8JtHzj3e8fN8yLfFBsQYKt3ZOZics284H4F40bs
3rWQ0rDXa85umh0ziYy3Zeu1AKRtZPEgUCxK8mxFf189GheTzO4juqKDBAlyYvAk
R+wVQpUpKM1W3lSdBNDaZC5Q+xz/4AZVDeRsFjm8CIJ4vAHqJJI1qBugVcTMjwnP
0hWU7N/cVWNzrCCJwqVY1n1Im6fdKyCTUcyq+xIE1LZMxnFyf/K2OxybxinIuzJz
E3bZl3GXFM8o0VInRkAlfg4Dw/ZUfy9nLsg5N7dS5h7jsMA6HYqGdRZw3RQqnyML
PtkrSPs83+WxZQCnoXFsVurkMuC14EZvRI5g3BtbXfuRe2FYvOp5DiL1C9ZR/Q4Y
pheP3bs/J14nW4372b6Hrtb5ny2/0a39vCNAnPTBzzDRuqDTJQc/0s8IFHT9EHlG
V/+w8U8c0bwexuzjsx+j/Gs8i/6elUokF9SFuNgTv56yc8xlcTOJT2qVWTZzoPUm
WyOmpByGsZniNN180GAJI0+/QOeHJ4MW8GBRGRigPBK/HG4CDX5uXTlg+7yTAZ1D
7V+lO45TT91K4GfPRpU/QAoFaI9GDbHmTjZuuZGJ1BSkNAJM/2wZBy1FZCpB9ajB
LmjvrPYBKHgAft4wn0R6c6T3/tmyHOnoBCH2fIkBChqHuhm+Q+t+UZYxfwlCMoNo
Ftsm7IAmx9teZkvdZy9DFNXo2WxJy31412EMJBhMdua4+O/Kd9C3ND0E1sLU7Q8c
2EL+jd4nKQ+zYlCoWsF9tv94iKw0D0MGDtERBXd447V+v8fNaa1w4PQO22Gr5WaE
5geO9DQoMgQpUOuHQy9v0rtsrIqXFiEaeXipGUtteAJK3xh8NO/EFu9PrYA63j9F
xgwWIM84QNnl1B6lgxSQHAVyIKgASTIQJ0QCB5gtZ1sS9xoolMJR0+bJPs8CMkb8
9V9QTu5S/TDts42nzVS79lOI9+ROZq+wJdbOGcXs57t8wmSef108EvMb2mGmfg5x
oQtCKDp+IPjZz/zbBVkdf1oQaqCURU6IwRF5yFm9dM/M0GD0O5MLU/u+kC861UkV
iiKnn0QdnrChXWlIBQ8bQb+X0EN9VxZdVughk6pLan/0hKV1C+/drqiGclNMM2Da
jEl5dzYpPKNBSe6wBfW07Ptxgfw22I+MLCwTaVbjC/i173KhyshiWSGjNpY8HMjo
V3MzcAQJy69oHuPlVY1dpRrbxNnmkGr5/nrz4lhmwUhQQPpmh6ETlpbQeVP2OU+P
PcMA0TYsi2N1SFqOlUetXfrbc8QwOBrKYnPbtMqzBBmflcjdIGek88l/q+mBcPIh
QYMXBW8b+xAjlVQf0XIjxWpzuCMHIWZqVWntwqlXUK0j4x9N+C3LxRsdBiSw18wI
2q3s9v/bQ8AL8OcKdRBgLm39CcMKgeXRNCcSeSDzcD3ohIS/skS8xB7Wnz9A/Ng6
8Pllj4j5btQZJDJaYnNooFDr8tTR9xH3WZZaJMaa1aKxgHdWW322Yk/vtcn5nUmE
7LnPG1WdJS2DG74zq+tI/NRJd/k0Me2unqeHWz5L41b8TTSvE8e0v3TVyO07pkL2
4LfgQElg5gBLAEaJYWRMVecsJXFRKM5RQRX+0tlzcqSUfpaORLUlfh6rV5vz7J1y
W/SuK3OtKdB8tU3cz1nyv6+K3AMRI9RMr6a22yuS+uYkjsDSW/nkzhUEYHUo5bsL
sMBRQ44W3BL4yhY1Z1yCqiPcHPyrNXC7ZUOZCPpH7HCCt6nJ9sYsfEEv7npP2pvH
P2vVzoRHtsxDTNe5bXhM32VB9+R3Gl5N2ArTL1brSzuz/1klrZEj7ROTV8eQ3DuS
irSYyQDE2v+Tc3N4ipvf3QiBUwRJYBxzrQZtUw6KVsPt8cKW5nkyyq5qBG8cLZ+i
UZHha7mBpE13ArtfNkwh7BkIX5xwZbFpb6qlZQvxgqNmMhG2B+tgq59C0/A8IWVe
SgBC9pA0aEuHXVns130itrda5FLCiTbAkkHY4A2vZtT7Lr6SKyHKbUxUp9wdn9WB
BWImvcyPjbnqg5xsIbEhz8deppBlzhl7R+J7zb0CElOhlP3vT+L5wDtO7J1czMm3
KMvRkM6E57sl/9RzCh38eUQQIhE+PLheOFy2H25p1mpuhlt4wGm3FvRVEpV53IT6
76yQhBpLcvKE8y9g0nGA9fyVncTgWzuf20c8CqyP0sYYnv1x8hIWx+qsrqjOxx6G
5OzW39b9FOjeREGI0nJIENJZy+6Ju9lFgRECSGUVAFlZOOAyDfrFJPf7234zI7uf
dhJXZSSzI4Y5qE8e+ojRpui8IZEKXRxwd0J3I8yKpSXMZoRYIq+NafwK3vp59wX4
d65PBO9fvyJ5dRoZEWj7PLo7CREyK4qIKNMzRoNau9GjMWhoa2UJSfOjiXZbi+fS
JpKH1Cr65mUJJN8zWmun9OVhMLRS8F2Q4N5FI5lRChr3/f16LcuCGKQDWOfTJSWx
81JX7bp3dZZbtRhgJYvQzalwCE4oeuvt1X/IC9S333ZOV7wA7lOMIsqzxmGbMVlu
BObTeRc+jJyLBMtHjUgRFVJnn2dWnKemtIhZGDsJxoqh/aT83z7QvKnfXio0qQ9K
iggWvBBAoTwt3ugMrsAJXUHLHm09VLNarzBkiSKC1JhKb4zR9mhTE75n5Yt4n3JZ
9YPmh1oVWN94b+x9qmT9rPpJTmY6LDGKoUJu7ORqxE0EPaUChvbPUeW9tdK24cG/
9TYgNAQRwkvuhe40JKfj3p5NONw/dj6FbP+QF6Y2nIsBBXhVcYQgky6U4V9rKa8Z
X7vaHAQCzFER9/P5lV5AKtf1tZQt0yyBpL2AsrAjpS5YUSVSxvIMtbaSONDFHr1Z
lX3A/Uek8FjEwsQuPIWLWRSLOHSUIfNPf3C1aAKlpzf7Iz/qG/0tgDPZa9V/syZO
owKN7qDzxKIdXp+AUV57VRrp6zDi1I+rIRSfAsftodWCi6takMz7nlzQ7El/pWC3
r6Cdnfu3FXCYNZ1+2A0yZ62gffqLiPGYOXEJfJXJDU/rQ7xLjZviO3R/4L/9MwKY
NswxGRE6g82WfsIOxArTqYAZ9XIE1ElWiRACeODEos5w7i5Y1/OZ8tnck+qvAb3W
AIL6OdOrj0HBaoFM2firVGcyIwlYerHG4ykkIFI9X805TUZjdyf07/1B1IsKctYP
WYcbs+FO9pukb+5IDAseuE6K4V85Sjv+HRTnI+4PqtGumDXmR3ZWYvj6Pbsf9kde
HOfysyE7GRudTV6s/Wohz10tQMvhMrNjQ00/u261lJUls5uOQBKd9IbAWUvIQKU0
of1Ri3eYPrtkFrmlNdnmJgRb1Iv5lwjN+s2i2rSLE/FG/kted065fR1/DapH4QuG
+R2p1nmFSNKG4wcWoQQ9CqitmF6li237UuHIx3ghCGciEuh9J1QAkUns0OrbgY4M
B9FLL44dmnQieeM9XgHlLNOj4BdL38ugoZQJlq2h3Bq0i90GePndKb8v/WQy18/w
zXw5bHwyE1zRb965MZtKT8vNfGT8dTbWu0ycs4Keiq2aTgdkJCefoBnJI4cRYIN5
y6ZnXJ16PQOYLHG9Ca7g2AFeRJkKTn+gEpZmIfU8yBAFr3qhxVWavTi0zGfWsnbl
ZNgDor6KFRk6/qRL7OKp/2SVD8kryEokCXHkhAXThOOWtkIwF0ql35qVNEK4zBT3
8BuUV93PYgHFWb9yeU0IAu0Zhleq154e6yIzjAdy8TrVlx+bscPozpAtWBo3pM5p
V8NmED63VWuLn5wBw1ier5g1Z6QBsW8mo/NrM2mqSsQW4JjSXubhiW5FE8A22UdF
semARugfQktPAWlLrtUy899ImoVt6BEpjsJjLY9DDqos6V6ABvk/KiZjHSGRGjzQ
CreJH1v3dGcYIbcUhoPCsU46Vzs23b4sF+7vTTo2kB4wEmSJs2U0Nd0MN5GQMeZ3
lsWnVDZTIi9Od3FZPNPL7RChJUOOIR71KBnkqKYYFx9CWyWorILch1bGX5KCF3NI
OnOIzblA1OFvmKZqCxZzSGY3WTyab0QgUYAiONkJsl+VwDCKvwTtP4UT7nAmJu2M
u5K2oIIjGcvYYrxDSK23yR40HcFaPSh/eXYZWR3EsYYRJal/Q4+a/0mdyLGhmAOm
n1FaR/X74m42UebnvKquMpO15CJhZBOYeuEHB26NlQ09TR151E/MyU+JsEnjpnHV
KA66kkQmcLb7cKQ2tsqrjK0iRLQxyblTMKs+n2OA23Q+aIKmPoG0rR5WNnbnBs/+
2TvGhs+1Cqhm4PLEUYzuDoeX0Vuf3Tme5LvWtlLtrQivW6+xdISF/tUl5oj7vof3
umINkIBrxDWLJ8Z/sNKpbrPbCQHPu4eCqB/02ZZAk2Bxs3uKyBqaNRz1qmFvpbye
uIpvC63ed5SESvu6vBk0nK3+JhG0xbXtrWEcePA3/OwC0nNQtmS+QrSTCJ2mWQhh
hCq/IfvWTsSPm/nCYsUYosQeUS6ZbocMkKkQeUKCmuR37zfdbDmiY7EGA2t7/v+R
uobVusErAO1pTOyHxwh/mX3EctUxmfClieVWIXK0B8ntAzuiJPWuhWyv9EaRd4ij
cqUnoUY6dPq12gpCf/NEmosx1SysP/j+l0pvgWZxWwc42KJfA7EwkW8O8RZgvr25
/rPQZtHe/HTI+RUEmFGs1TetLP9J8VigcENdQagUymQ8nf295Ic+3EhckgGVbM81
D7q4pcHTynrvOZPZ8jDhWQpxyf//ky5vBfXZv3nkvdHDBfXGH5JM/RNX0nwN9jGi
pSOwBlMBWz2LqXCA9iD9l4YEx6C3pYX6bpRQaMMrDndcUQMnSA8FY8XuYRKuViwm
U9ECHDO4mfXnn+GRpR6GLdSswt+Y+7d+7RypXxppPRcFnKa7gt5N8ebiLkC+q1Li
GrDGWZYjhoOtKpvFzgx7U56Jb11zH+9XxgV459qxm3/gq2Zd1jOSqoRxG1Hdr+F8
0OuFoJGoVvyoTq0DIUncxfeK/CW/vxdY2FXfY/p3r5SCZG7wn3MA4pVLEzjC3C7L
Ye8xJk772VpZPTd5pabEvJrSpGhq82knYc/4kfBaEFwZXNZEmWcvsYtjSh6IDoR3
LF4U51E1WA2PbOmIb6rXtXXHf+vWlTwN141IqOj9MmjDhiXXmGfQ+BB6lanj/Vuz
lu8Gi955F6ERU7vQjozf0bqLNoMv4UEXAhKW23Ch5ILNyhTyhNR+pzv7oZ1q8/vb
8fOs0evsNVkUSkomUvNZXrnW22QwTnX3OLHu97eqdDo1xMRANSovEigBpK9sp5o5
SVo5N7+y0PhaJznPwD4O+7WN3NWTHuMhgsv1wYqLFFZsUjelqScCRgpD3cP1JDEw
XfPgekrym99gzcWd3dE4xXCVlzV8eP2Z1nuQ4Bk9qM9s3O9dewoE6zvaY5Y4HOhK
B2mbZCfnFdpfdysy63apFLF1+rJmhgkxI7IxqRqILsWSJnZMZH0HdczOh/jaW88G
9Ma5nnjvmVyc4Nx2fISBYIUDxIeE6jDl9HEwY59eDmJcXEzCxCQgjlDrX3akHQzd
lDiPj8mgbNj1XWrDxFTSpMJYRKMwjiOpO1zRAnwoWVGMfqZ/vqHSHukFrJO21weO
LjIUZ8HKT0SE5dUotDgPuGFmIV7hRGZ2RGe3s9NcsjLrdQjtDNLoSrSRNAzF3Le9
ShS9/UVw9FPl7Dslcd0+GVpyOYSFLtQZvuhzc8HGMeP04Mm4/3H2q5g3FVHn1ku5
zEb70LyUvrEsnQu0TdDQ1qTjSvIDwSavTP+XsfYjbr+Co6fKOXxCMsCQ5dVLtmw0
euF5EJWNBV1ODHQyU4kW+2xJjXRkB6s1K/9D2CxUb4Mf/pE07EvxIIvCoMz15nqK
AdW/zKZaeRBeUObGw9u6XDg284WZ+qXT1P+yLAGS2EKgkqviafEYwICNhLDPX8Zg
XclJ6d6JfGGcMnG+LgJ+ulL1lGMYQd9Lvnx0T0tXKObMCICGBaZpcUetGO+yPHd2
VOccdGIbB0lJdT9T/he4LIaKNGHmxviI+rm+OBIFOQVBDlQ2VNMVb2dMH4rTKgab
Gv4egyVSPG7/SE6n2/kZ8cxn6pN1V/0PQ8AgZFVSgALGxygTURyD39fKuWdcytsR
oiBMI1z7zsCpknRAcFR0gCJikKuf/vr9zVlJwuNpP4sx+nMzvwGa8Jz8a46JPRDt
hJY0l7tThWjpVzMRlFbcbwtguwFcCSGD4HiY1r331aX4PTi7q7U3mkbkQowz/ugd
oiH/hPicvd8tH9JYRfwX9IzfZj+pjrExmhRC8mjKo44aoZJ8cp9YvuxVjKi3vhji
dKn0bsjLItVOpMt34xaSpHenmxx+T0c8My3ZVDwxzh8Q7xhXT2zto0Jf5V+F2mCE
iBfswz2EAXzLWPrQBERY08ZYWA/wdUuIZ+LLbHuSQIbXh7COx3fAxm0RL660fiEd
7WaARo0YJYhMDSOyYNYnubZcQsGAQ5/mDJWsXPu2o5Uaa3+Zl4aIjsM2CiYR2yrr
HCapq65GKe4qwyIFJp9207uWeHNiXSnahRXsv+q4wc7s5/HhD2AuuEFleBYrEUQL
YckJ1x9zMkA7T58dZFTAy1Jp5Ca3d83r1GxkI0PZk0u5I8J2SnwISKGT4TjzbHzX
0EyTRgPyqyB9229U1iw0iqSCHPFXULiYWgMCcU19g6+WH//v4HyYEAvvQMwtQ28D
hF/amOFcgm59J/oEHMxNVV8mzS3G4y6XI3NWsemKDeYfCQK4dkRQjTV6mv5CdRDR
zHuFBw+yE6ZTSqu6ji1I2G6FkBTvqGg4Dp6evsnjVljwiNXm98JY1g1Fa4/AsEWA
X2kNku9Z3AS747MKec8trjPZ/WbFj0CbYa42MIf+DBrxWkHqaaZhhpKl3sotGZmN
lVUGU8gDkSKD9XdmeuhUyI4iejJlNpicc30GOxLQz+YinU3F2aR12dEDNOsU6W7f
9+8tmerMqMFdm/136QgQGKi3uBPCdh18knuO1ovqXQlHekhcAp4GI6s8u6rpqEe4
1eUculXoBlx/EWda8y2rye3IcCiwflkRtAQ7+I5nTsEMVHhQbmkgJu7mRU0IE9jn
`protect END_PROTECTED
