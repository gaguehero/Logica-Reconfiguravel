`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJiUqmxZp3wViQaDkdo+mLBHwNtSA0DW4XveNRfffc+yt/gFydEyWK/QcYpY9rSC
JwQ6dXHKFmocKnm6Pwk4m4okn45dKr/pPVHXzzPqn7YbXAh5XExUJMVyE9UOBi0y
fzr/GA6BGpRgQuPywIA29oWVvVVwBtV7rzGLBGTcsYMmrz0RFKevouJK8Or1fKnR
+ZW6Riua3EJT/aSrjXivJHdIjo8DgKc+FH20ORm/r/OVhonMbR5JkuGGQCcjvzBv
MLIJRj8rOFS9ju3wRGpKmX2ExKi8Nf/aH/hWIBHu8Mpzdlw7KPnFQwFSIBA1s1OT
eQ84sPWIRm6s+/3rTRxaS0Rfd2CjE/g6m2AQsnhQZmSU7aUKjZAqxlQ3iYLsA945
bIagVBjmAk4ywPml83rtUwPVr+Ssrvtxmj60j02W/cx1sJunkiR3kib7zJK2mDyo
ZsSQvhU6h1msRxY891JdDIY8AaljNKjZlls/YV/1jgTiw4gdU7huwwCZJ5cBv9AW
VIB47eyMagMzvB5R2feOCgjW1sCxaTATYd9ccX292VMM/cmk3TMpxgDeiH0wkBW9
VEaLySjRH0ln9MNOXtgqjzppznNjAubY9DU2wuTNpULqhmPwIR+Fk2C37wKKgR9S
hSHPcJahegImfBkUniHx8Q0lTTomgllkptlX+EZgxAMNMBtcDApY7a37YanarD1N
gfySSOZQ0+MYkZlCmjkuSCCHewz4CYzMcouHxqvT01IXSmwRhizmm5mFf3Ir0LUe
y2O6j5a1s08h8ZdWLuA+JP/ktEC382vLJNqiDUJpij2r4lmcPqXp7kIY5OvHZvVz
ZDUuH4zyLZQVG21/T0+k8ojo8Z7jyFGzlDs/E2d3DFilcrMnKN3W8k7PHd94ctSk
NloLwiarcCIMKglUKkidzzEc8btoSKMDzkUbkY186av90IbSemGSHGhYEeb8es2j
nVoHglz/dJmZvbd6XpxkiBGyi+Vr0ah3qmPVj10x3iNw916NzSLveglafNyskzbB
uy1zNg3O8YMtpYmb3aKzcbMmkUdxH9lkMK04/QnMOcumr0hkGVY5yIi81qtLH1rM
VRVzmcC0EjDGe9vpIylIzjTSs5eXIrQCbDyfgjsgPklNSyt4fLXRqtg6Wliniu2r
e94TYyCPKUzuVTEZHNieXsOxuf9e3P17xkBQfkASWDnET6RAJ0hKjiUSaD4Ud79z
3D2cCto3nZuRYHMesVAbKfVUZtVP7fmRqxqqWcznVfNGspVr8HvzmDA8h5vRmfu1
M5ntcLJVSRmWFTsBV5YjWGAVrUv8JDu4RhyEbxU8E02ZhaQZeSegaIGWG5urjGsg
emUquYjlnqfr74c1eLdYVK3cdTvccj0a2hkQwimVLOSTKT3ulIZWU8t0aQsvDtxD
nH75V5b+u6Sray23XlN6DQlABbMsTuY3grmw+NuYLgLZoPRyozGSxpn98unbp3Qx
fyM9VMDP4wavbFdv7iWPa7v9son3+0KwLaaOsimLz+F5NMBPDKbCqi6nSWQAVdVc
Do0N3FiPkHM4c24Wp4J62Kq453gjWI5E45GbqErxNiwkQS4tLF7ks/t44JXwWWci
TA3c0fzYPBUqsEPc+n595QFRg08ST3xSHFMHLspzn2S71Pe/iDPOOPNw6A+sjHht
oDiRhh2dVTySEctscpVv3ajMx2l2Z4WHAqpQ/Ebr+ekOidjHwJwwPJ2wIXn4zb1k
KBx5y22whkJrGuHvngsqLV1Fq3d7c/xJzfsekUCDsmFqF9kHpzDCCL4zFv+nxmvP
NFKR1OG9YMjxnLg92knu6g5zrwoNqi6PDlfNn237cfnzsa7HRogj+goztshEqoVn
5i9ZuZxV9IvGUL1RYjoet1mPFg3OZkfsy/Hbd1wvGSASpIQICA7NykXStAIMqNA6
Jrh+j0DCHVTumXZ+QXEpPXVgyQh09C18ogGTsyohJEwfiLaJ1madnjdAUK9KjeFL
IPjZCQJy4RCxohZnMR5rFElC1cHMq8/Q8ar9zbsLX7yml3nrbQc9KcLLojZFMPKN
m0pDzTYjnJns4XBulJu54mJ5J9zzIw1+Fo8tZhWtd8+JdrzY7dU5iVRBlkgDxdVR
u2g/x6PwApJAN5Iri7QCSyd4Tb+7/1r7Q+bPioxviHIzjMxTJbnFyG6Vo7ssn7NE
OAzU8cRdHerYIdjBQyJalYk4oW1mczeB3X3gVzVwGO0Pl7h9xJq81qjFZ4udV5QK
WBjIDzSSRjqb/jN0icdIVpiPEWVdfsu95kkR5ICHt337oaKaPBtBMBwVSZRMEoLD
4pYnWYGOiCgI3Uy26z90maXYkFeL0vTWJ2Cob3rWvNd6LAKk77RTnC8aR2A4joiF
Q0scp0Lm8C4TSiyKOqjCmrFVh4TH9adxT76EPNyhJMp6rB8dVfGkntMuTV55d7Wf
5+8lGWnnmAnLL3oJJG8axJFC1Q63HgBPJlnjBr9KoOf6VuIW2IGV/MzuapePIzN9
HMD4BWidcnTLPPM8km9RjSKIWpYXUvt7cWD1icwBvvYdBw0H3I1nOLgntHRnApCC
VuyqKbjab0K+EqB27a21RXpOqBMIHWDZGFY7GBulnp1PvoWSrhfqIpGrKoVU1xpC
dpHrTR5DP2xdAXb+Qdr3x0j47vNfWQ3NR5p+fpRNdEcvODUbVEu7V2YftIfIMf+L
erjEfvDZ8f3JL+Ukvt0kZIesb1tkvZC73sbL0KK8y3CJvHApqc1r0TE3iDMSamoD
3qsEFnqjOEc2droAehz4r3KETUtilLf27vvEC1w6HyvzsW1IhXTJx4RXYJiAduEy
VnY9t3hM0oqGK2KyUGfdVd2fnjjRIDUnInUddci47xME2OX2yiy41W8MRxrLD/MA
kOxjXM6GLs3zfK79zJ6LAZw68CEIVMz62ySMXcGRQE7jqe5ckfgSbfVz8GaP3qui
Hqqx6LilTmmt3qGhxNYx7VHEGgdOVCigQCWTRhZlvgZNNx+ehROF7VdUMhQPIdv7
DwVZyCDHwv96DQ88XLkLDpfMN4eGPhc1qB/bpGmldGFvQm2vBgP0hvmC+X4lDilj
8fhi+Ig556xKAcoiedCoAtZzu5JkXLogcEQmi88Ibkhea9tZ8tF8x0yL8IX+qdbH
csA3IsN618UvJOYZVa4N2Cp3A2sA1TaVj+axhvnuYNwQGwwtJcgMBW5z3zSzfTyE
rCtDugID2vlnFOCtzcMq4ZIQZi9khRALHrfv5KxzVY+yVSfdCvoP0aVpf1McizKE
dR96NbszSx3iFIWkkVY6Y/07P1LWUy7LbZUgIcxosX/x5nyqRc+4WvFXBd1gsMkc
/8N6Cg9G0w4yEtUdBPa4DyXXVslJ+bzwLSoRMxGmXNgqkYrvORcCKZyZWRiRIQ5G
LXY2ykzo8pxK0HHoyyEzH92Zr7AHdgM2xMW8PnYfxBM9tdrqR2VHHIc/v/wTe+nq
xKzlpVa0LHQ7VZqEJxtKRUHAHGBxdjTcEzLou+nGFX/4l0X2KyMDY0lhtAl28oIl
9ei6rhdQDY4lO4esy1qzs3b+u1P433pkyPC1pDVCmEoQBEHKEAQ2NHERjj8095Bk
TgB7+Of7sPtfCdEPYXFIHB1dr0iQwpi2tCdeTWZlkXVDH9IIJviCyOAhkiB74IaN
hB5ypPGlG4ioaJg5tBt1//677agoqC1771clZYbFjjDncXg6h1HJb+wV5yWMkcD0
D43shfmcaoUTN5Z5zAuKWm62DCuGgRI9eBPN5tqegB2n/xcbOSJXN4bP88zALrsJ
Q042n7JUdM9aXkqD4T821IoEfl55iPUwLQTt5lGTVdX2WxYo+5HQPZJ9/lIWdZC0
zK4foGg33eVs8Ii7mvQDhCarg62NlyhEaarhqg3VpNuGR47qaPx1+XUBHh9FTDvb
zcUnlDPm5q0C4IHnJrpjTW+tzgVGrg+mv6MGORz/pZiU5g2ycOcU3HoSP1E4oDKO
CUoA3D+++wkjYudjmIMZuFLD3DL+bA1svOJZ/7xGEDfmBINhsNVpnZcWQ7IK5P6q
Wjqszs8R319cT2Ow+E0R3t7MHhba2dH1RBckkrFlj3ZNbSuQTHyeFIk50F8ImjSg
mEZESKKHI2MOwx0biqFho5yvWSfa0DkowtDk7gclDH+cRNhbEX6veF0rrgLOij6M
fI+C4pjQ87r/hMega0fKxRnhvnKw7/ZfMAwRLaR5DrW7ZilXgCCiLotzFPiSrCVX
3X3BGD3B+fC0MgNNSUZQ45JljcPmnG5GvXNU2SD5PDtjx3TinLMp1m3k4onNt4ra
76y27VQkRsxX3IuvGXvmPQI1tnBoXAzRplOJCBMz1QyXW+G03BZ5zfatNiFrsyPF
XnSE2UfKChDI1y8UsO1yDwcX86YmAwAEckNp5onqD/6xYlYM8Mn9eXdhyqkm/B4i
XLpfqQbXnPSnk79lvw1J+KFWvDp/T8OQn9+0VIhUrCVcDP1MR1A1azw+lDT7ZMnV
yxyBdSo1qMMQSeV75eA5/YNl/Fl2a2FvOggxgZ3tzLZ4wxu+fTEVO9gXMI+WYSqd
7A69CMSJHyEc0c1BEE9K+dzZF48+EPd4DEo0rfvy1CbG4hl/ifvjxiZF7LKKWk0m
7TygAScpNk+49XXSH8dxLRvRiFH0R+czZmASSfZnOI9IQV4nOeYsI2z2WDeWlkZa
+sM7s21a3cMBUWDePjFpEss11hNIWa/Os7J7FJbyZ9AEmeIgszSFLq6UNWJ6ACwm
t2VwrkS+D/aw0inAFadhSKRmRHPhqF+taYd6jCgphtDTGD0XbrTTW7/3s33sHTOc
ZavoAb4ZltrnGqtWJcCx5LLDafya73rw9LWgt6c/1hyPAPZ5zu5j7p+3OwLJFky5
lRuHie9xyinQ4hrFnj9y4hzsWJREDPQMScskKzpgkDa3sSgbwLlHp2TP/w8bsbwk
YZUgDhQkxioTv1O7lTixx7lbLmDM9+cJ07scj3RzYXdaw0PghcERawP4pjQ3eOWr
57aovkj5tIvMzkVN4pCcY2C94tQCC6Hs/fuSyqM0EyTyPvutaKLJNt4Fsgbmy3p8
/qQVIt9QtS86ONoqwP0k6/izm3jJyJzc6yjJWJhO78fsYrX11nsD4s+2FUcCRv9w
w8Bxuohv/EoCX8p54DbKnmbjDHY3iJn3EB4mAMGSR300eG7CyW41slzgv+LRDhP0
IjYdoAK5HPummr1eeh0x9crd3LZHkSUWLdoOZqc2Rs5fa0J4L3fIEiMiP/cQmzPR
wUYZMc+SDqJoeK/5uvql6fWg1DoofKeY+NP8beWJC4EVFDdyTiyD36VzJUV8RGic
qCN5W87gWxhxM5duyuOXWIDMTJW2fxkP0JjTw6s8pu0EpJNKgYzAuo+8WUYM0Egd
Q4XAPbe+ZY4W6psfKLfVPKoiXY179Xibg51LEFa6PfetBnPsKjPuKiQ4IiMknRnC
7ZfRek3999aK+oGMiDF34A+NVwUCHE2JZwqrLfqdFp7uuXkmXmXmjDhB6dGrVO0n
dULmbu69/aiW7jGXfAQGQ/qfRVrWXn/M0kbLThPdmh1Z2hRR6KeuodQTAtYTDgwE
xXsVBcWX57bf8bAAmq0DmyPnsnce3kbR6FIZcgT3R0df4cLjHHG1VN2ehvFZOq+B
vETwdPe3AoMtjOUMPHYoepkOwlDCXGjnrVQy0z6WHmpRBVaY7J3U9UgjJNLkrccJ
ioLOR1cxPs87MOGZ6FnIqtCci8SYuHYXvDyWGYupWgMTkFGSpAc/JCzx1iYArHcj
B4BlkmKTBPzRGtPlNrOP/e8dqW4JjJzTlN/aH9JN+w+F4n1eo9St3mrKiKWO/kJK
GLsm3pyAjxbFyMce+MPaLw2hRaeAkL+Tr5VKrBjyjM0U8K/Hn+oiDGZ6p+fLW6eV
3DnW3Ef8vh7eQzOZdTjNT6LiTj3+Eue5LpxNL3gV5O15jD3Jqzf0BJpzUkoQ7z5a
aMcmwj3LI0Iq/upacZryrm0Y7hScNIo9an2edFdc4pbzMSHkgPfgq0iSBuKhHQsW
vq25irYkm/I1ytp8wMEoUo7Qxya4tw+0pd4JMv0pN3rGzzh/PEKiSFelGc6C+b48
USqrzYtRFSvNig5ZCUyOTSHfP9GYqbOCxpHygaQDQboMpcCJsn+JjlkOH0puARM4
vS/MgZ9tkMfyICLVwzKqhk+h4zm14mP+bgmYIFDfW/7s8AVir0UMOq9Js6XaUIt7
MFW3B0aKtRkYglkIMiV0UaisiaPU3uoVoS0lvykBu1unyAfdPQIXfy5M2BgVSesT
/1JNc5o8NtPCHheQQouCw83FnWNk0dlsG299vtoSLShxwlqqD+WRvo00dfgPN/2k
7nbWlduPueHuAab3e4DDgXfm4Dt2CGDrmf1BEWyxGxItTc+6I15MLHqDbBEEl22w
ktLoquiV7l8iA2uFpjzbTQkicWBfAjAAU3AXeDM4IXhScQ0wEfNFPR8W4nlxo1qG
jIuWya4Dge+UE2nsbst2g8oDSrTwU7otFOXcf+H8UE0Ij4V0snLKI7d1UTuNESVT
SUp81/+axZdmVIke6E2GNN9LskA01vGbPFX6D5GLrO3/k/82hCQmh21+6tCnI9JZ
9js5XwW5ugd9lQr6UdfiLwGOitNprD+sWoTHWxiFJLXOTwb9BnTmcNPuAq82Z+wZ
gkOaUXa41uowTF1UzXDbwIikFAjQ6Qb2/mkLdMANZT0=
`protect END_PROTECTED
