`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYazjiaZngudfCjWj4LNCHN8TpjHtzQN3KS4qizoetu6iftKvBcjtpW3v0E2u9Sb
592QNKNM+/rZ1HlYtphwF7N/gFFWOb/Pr32HrYHMe6+Pw/A5RBdYv9NyxSGKfAO4
ggSzpj3E7ZYwf7P/BmxyA/GFmcMRgRryyvz7nZ7EHo5fbibrAKOrHNmPXKUIcDNf
S18xvP8qEc3O54dRNzAqQC5kCrnnZ/TTODxqUy0kLZ/LX/wSEFqlHYWhX7Y6SaDw
oDcNJ6QZb3VnA1/QurSUqcyQPcDP+ufpniwTwAF4i150t+Se4KGNXWsGz+pt3qnu
6acG3SFSXIA5ieHraYtTbt8fEnVPiyukpY4FK1DHH/JKh16IH/vOz+Cb8dkHegYy
R4xyMcZbAEUXbx2mT+t/gKhsUoChOb19ZcWQ2T4B96UQNxg5JpeihY5YqtyhPApe
MOqNffMdth+wsuX6OkRAFB/CXTj1EDdwSV0JAqsvuT4I9jNEMlEvXlIoWNvvHKAz
rykN38MPHlnJmUTOxQ0CaULrIjRojqmbSEp0+Qdstsp0O4e+oVhfm8pjS02fnG/Y
yln4dtLGGbovNdnNS3MNX4EgTPREZcHAfotYfUhyCFI3zodulR79IsmfEjGppf7H
W+O/+FFfAjuE3Oft7UT81EMNIDTc0XBQb4q2+ByWW9k7elLve5/Oe1+OCVRE5sB9
fZMCDnyUPg4QyZF62SOvjrfTSYCcghhI79nQr9sVkP2laxANk2P/OrV5qh/meiUD
vpivamzektKFgaAeXlCrAbph8xu5gQh890t1oqXd+EpjB5oNYs2aZVzT2f/UcjnE
CvaFrv90FQ2bzgxhIOIg6J05m11ZTZGWB3RQ8fwKm0dUkwOHRRzoLHiST2mpx45W
nbRKkcygG7T/Uk1WQenxHkHJV6I0VtELDGfxJb7PNZBxgkyj2pM/gzlur7wSe02y
AlYRtWD4SNs8ddCPs79HCwL0YB1wZuuV3gqkcsXFRggHwsFNBeYjMwAUu9ihvi1H
AkT9V/DADtD8RztxdTR7kk772OM3tOzXHrQtjf9Sc8GzvBoRKzQF4F+TMaMqCOlV
1WIUkejLhBlrJNHuhdKVo7tISOQsx7IoeI5pLMC8JyeuL+XHIlWZ/PbJkAxEGi/p
M4r0XXlm3nj81YqIQmLJWsfgXEGUdS6Z6hSrmU9bx8vFwmpO0aMR9ejIs2IF3sdo
zWhB2Ps3AwDxzXAZJtIZNKuHNFwMqAqpVrjZPVbmAmahJQc2MHcMFzL6UeVpqed+
jW5Onh+kgSViQlxFhO6Z09pm2eo1HKjPBXFw161FukTtLUCKwrba2f1rhExe27Bv
3kdXuMRAiLL0nyj3WzFswBaZK048bEnYyZnes3Ls39KoD5feZ3PJRGjq1G+LUbdf
LM/RyGeJK8Iuopk/S1tDog8uMrrPmnvjks/GFStAsv2HRNKT11X2g1DnIiZ39BYe
X83ZBfgXkf3G/nMHjUWx7G2iQuj/4z0no45lHMtL9i70JqqpO1kg+RkYDAHdoUZd
4GSMTdvKRCGIX/Pl2xJ207TPKOFmBa9mSljuE7E0zz1LZ/+Dpp96Y5LE+vOlN7xY
Tm1HRACGscl//0RPFYp7g3bXTLzkr2tFMm0GbKC/zElzrCymIKzBJgLNoKiPPp3B
cs4GFqLWYS0F74vrtfFRbb7FjgHzI1f0gajUC7D3NlWAFbXRe7IukbTA6iK4tt+2
DugXaG0xZ36AQI94XHfOwsoaJnr2IRuDN/V8Gj7L8uNmgkuIHOycrhwkmwGsHx/I
nAbhaKnpRBzrsffq9sz/0FSU8fkGMhZacAAPB/zYFw6y6wNZs7+Wr1a/J95ernHc
YbFCOzD8mXAF8Cr1h2VScUMuvc3zttfYP4i+/L+8WRBWF6lH5ZO324RQATKxGObZ
Kq2t6YumlBSDt0mmgflI3SgjGTU41fDaeW8TXHRs+AtEyrq1fBlSJyeee3m7PXD/
gFZ9x+pQ8mWYvkrvDqIemxD3l0l1Cr7N2RZFsHZ8rxn+mdAEHdzlecd9pgn9LEdv
vWW3vowr90pU9pN/VXIU9Toajpde3Ucait+4PT3ya1Q8oBn/+ivw5PCl6kP9NxS2
vG/WGrIfrTX88wB8Je/9DVQ2eLwi3s4mtc895Qol+0imjGTy28p8mzBblyE9T1Gv
uo6J0ZuZ+MkwAQqGvd/flaoNev/FvwZh28znP1swKlKKtNe96Gr9ONMjYomD0Yas
RvDIPRURze0XXr/s3iM4Fg==
`protect END_PROTECTED
