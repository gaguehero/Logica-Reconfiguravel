`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMEHFD4grrjCX1SYkZ6NfJlwvHkfBTX/xiP0EXmYpox7gMSSqRjgVKZH5h4vN0a1
FJTMhCDi1peztIIip0axA31iacz84SkZpcPdzWm3PSFKQARjAWSYKZtQWI1kAKO+
oSOB00zQx4EY1F626fU9Iihk1Gqo9JBjGWlgf46uOoUiQypFNi+cRswzyP9bVF8e
pW6YpvebzQTmJIAduhgbQal++zZ/R1HwUSTuVPgXzXrxXiD/cQwLCeAAGe4VTube
6K3Ra+MwzoleZOsrcgQPUEtP94B8058MhdGlLW0FSG4va6txh1rxUexsKr2qiqG+
IaZ8a96yZllAniyjJMUg2l8hpDSum5aj9rBfNyQTaGmR1C1YqBsDoopj/tr0tf6f
nUoarXfia5xkC2SX/Gbq+fPTdujP2i3MsFP6BjtBXSoiS+qCkyswJ53YKb0z1HyH
NFLkRTWGZEazYP8eW8bHGwnDcrQMXK1qz0VPR7+xWLojEEvnq3jZnIg9Lkw7eBNt
WElQQA3Mt48THTGGMTTcmbthisPUkMfmx8bzk5zuoWHeSJRzyXCUrOuKDNp0l/hi
2cshMr3PnVlNGvtT4lBFXsegwFwEo+YnrN2mfB0xqi6yHZZ8EGS9308eAq5BwLu9
E15zbxlhnmjAkfAfifKQ0YSOOlfhQHCPzodmXIyqQmp9iNffMFXVx/vO0PqocCcv
9UmWB2kQFRsff9oHPLG5yD5WQ1rOb5CeYaiRL5wv49A/+qCdfWfpmIVeiJaxSoxS
8/vuD1baVWE8FKbXkjRU+uIxUxlixR95h9WmznUPD+bIsT3LBa2XsIFB77e6wa3p
LdBnkSfQb+diTjoIMWsAOmfR1NTz+3231wL/UvfRn1bpFCM/hrhftoeyZfMnso56
1rfsRABRF1UqGW974vvqP+0cCbbkjYymh48SnPgjz1LsD1CsPuKiTG/HXNusv5Xw
ahJVV6WVNH5exBHlTookiCZKIvh9NyGqjtgl8IG1cNoa+JMUsmK22m7RxMBVeSx0
3KSGD+Ct98JocMI2fzKoVbhQc5s6v8vsnDzUbZ9OVBjDOec7R9gyduTZFkHO8OiX
TvOZcT1bBAywVmYwXklHDffJSuFBwoU1MA8Go94dSZ0uDUawOq8sjOKJP0r58Dhd
eKeoNUUy67zsyA/Nh1i7L5JoI34nrI6SKWagOwuOO6EVTXDbJNJQCDXjbYQzpAe7
jH31RxZA4mYYCVPboGSFZaCE4qOWvhtSiAiiAyEbOsW4kMKwx7EmPlj8zRI4H4T+
OCoYmeGWQVH8gSnBG9BPFFw9Acphgk8GT9TlenKvL0+ZRHf7Izqfi11vnmt6CxiZ
rf+F/QghN2LtkXWC49MJReHIGcJzm0fiVXBR/P4siVix+Y8xfB5C1EDZOKhpC24f
7PhDF6cQJMbNVWj1FSUtSja3xLwJ/RTSogyqRiSut2fOyvQ+B1/7M5Sf5dSJTR+1
F05DWxmukYDdeF24kFCmQZ+7i8oYDR+CL/TLnTP/WzK/6Z58GBqwMFG7OmD2WV8L
PSQ2sl2CZabi6LI6AEzkKkzSpvI+DrLO0LSg1rA/pGT6wENhESY5W94QDizyzlPK
UBU7vByh01CWZ5o2lr7K8Kiz3bJoE5uIidEW+taLLVLLigI30KlAALHLuRfAfg0g
DYxkED2/+Ew/UUkDLn/oaLZSM+25TotLmejD+RD87GlyE17CCrMEVPor40ESFddl
wNLZqXXZT+s6qy6bmzmTLgNQewDQNhOS2NbSD5HoOr1wQBJhSWM2PcCpggEMjuC4
aaETOGhKwQ3aXBYkHxJEgTfhcv6ApkZe2F5asNAmu6AziT8JZOwKhxukjzZiQMlY
4VgikwrdhScr5Wl2A8qebm/n5B257AmWFA92JpgGiGGMKlsNM5IhmT4+Slu+XsfY
sZji5JpKxPKLMue7YfwGi/omwywDrCKxlG6eJWRQIKY3orosZq1YfLh45HRCXxtL
TJ+jhCyACM1pYzxSzHkYMzwUqB2O06MVYY2iZHUBo61biYK/Izl5P825LAFKClGr
BKkFVqMBiTXdhwSCKT00afAqNdmJOFy6VekbUvigeXhThVcGqsdM41wDUUVjmXvr
RMGz4KfPDUbbYypVRgnUzVBvuQk5rUcvBqhlCAwaw9DBETW7eq/mvKOomO+ppwW/
/79eohr1uPUgNdNLH1Cl1zu/lJ4hrT+Z2rhvEilrWq/wWcCc/g6AarzSDPaLB5rh
XPj22K/YdlJv4otwAhKbdaXEGTidbMNevqwRBdfcsZYz9VrzYBxqeACd1wVNaYRC
77MMYwUhzt5dM5VLwl8y7O4p1j1q2xZGBI6TaXVjK6Oo4cf/o1yVdbDKIvfmLsQA
zUy98YWY0PeIVo10qSSLd8RvdEeMUTdHerg8h8GVclX2GLsw/EDIWPw6HuKo+mLC
wtX7wCYPVkuTVUiiTBD2xUbJtxAsRiU0gzd96gtHwnxSIvBtdS//hEvzOmBVODSg
GByA3EsicMD8JANYT2t/s0EsF2HfH2/kRQQ5y9zmOJMQdOKDYtDKItfEPDioiKrp
HLs+dTM8Hm5nu0n9fDC84Mje9+J0EEUSaeCTHSsWvaEWPBOv1g5Z82tqmJ8wNRLH
XvNRQbiptF/AaA18CxJZqvORDd8ElPoAuUtXPzvdDADkcII0fPwNwtPbwjLEB/Ja
cwim2frd4/xbfrkMjJjfJ578D5kyvP+s8ePLXCkpn6XJYyK8vYAAKVf7NMSCfpJW
eFP59raQZK1XiAH0zb+d9h9dZZVxy49sjVfi2lyVLZOb+qnCyuhnZH+a62fBAQIW
n8Pf5yoPiVvuUeNpCrxt4Ph/bvrmj/bpZX5zxsB4jcWOaRuzcO/p86ghpvHzqaaE
GhWvBAeoQGIEFGdRIXp9Zph4X/9U1bmIqWjVI+CATl7MipvQkn2iK5Dq1z3nOJRc
eZi5oaQF2Of3ajpoe7x6iSNXycGKSYwexDBMTUtb6gsGSLTgvFOBbPPuSm35Irsl
HwiW57ucf6y3zG0c59B8wGB52ZZX1QXLGUzI1JcCDRAOod5Ad2ladsyGRKdbX29A
0u+/6mrkZWqhdYDtJ/Szoo/Gp/d1qIAMDEYnjmRaEgvQnD4gblTwTRklR5aNraqc
LJh92uBiJNlB4GjhQZRD7Rg4REVPdx+Wpf5nPMLe1MlNs3Hmcszh961zFpgPcW7c
Bfc0Ud7qx75O2/bfxrhjYXTZTO5aUxeuBpFYhtw6e63NIeUxfwaH+5CF9qWguj7A
l64UFhgZqJZ5uTwQbZ0SfH1DaUghpghrba1KN9O9anGw/vlECacrE1ejN5O3wfAv
vxkCIidijg8FBqffpMHdm6pyXNTBVBfxV8dHTdQRYIhNq9toH20EgiAQ8QVZH4Kn
N+tLxADXeWSl0bbsRP+qg8DWQC+1iSjwpsLKdmYWYk4/NPs3A6jDMGFIqnNYeXtQ
6DGWnyvAUUVKDF8vcx5blTBQBJbvxy4U8DPneRqx75QCLOfimsf98jEWceLTv9hR
G1NmOUH69U6FzJQum+xyJI+vEbIMSYAcPP9HUIvDksMaWJg2jBWaAc6mDffrh+xw
c79XNIdEvgbyj9V29SzU4onCHcig+/ud5GibwrI1npEWLnAW0r3+3O1XwyTeT2Dh
f9nXI6F9JxUSaZqKInw9yDqfMikcNKx2j6AAPIwIAwHyvWRWUJwp1HT/EzB8e/vP
IK2U4cUnqIqDYCRKFvbpXbdV4aJyVBeiTvePJLhPCbI2bizT/auCgBVMLDaHj7K5
2d4xjN4u1ItiNtjxiUtlv/cqwEC3m+VPpyOcDyBpMzh+axvueGCqAAUyd5/rfzAr
7DlqLcedaN2LrWG7BAwOqmxoJdSOt8ddijV5hb4H80mI5uIwnU+zV+stl33GZgvz
biKQN3Uz6VkUgSKASp9VSPkt4aSuCtUvoY9urv7Xj1eNv/tygmWzuiVWGtPxLg/f
ur79yMA+MjMk7p25AorxJjOQJp1aRjKmkoJMYn1Qv0W6v1tJhIGHLXNqreRIdQQA
zRrwO8V9Fmm0S0Cx4jFpT6msTbRpH2BF7EHc2OD8NlSkip8YZ/LAtXBtAfPHqapr
buNKASXU3SqrTG6HCAVdxAMb4wJMsmr42q05gRQNAvyFV6aHQVnvG5+vZ3v5rMm4
ApxU3Tf19UjySYyvPXU2e2aUULpyM6U/TkxSywQj4akA+lWCm4e2RKnNLsa/J0L+
B8gf0q/GVUBpaeXZw8KfElAflb7AG5B+aFal9E54KXfRhOWTf67FP3c/9DYDBxhK
TNK0A577x1d5TvxAMzLi+1p+G8TJLtCy2ZehE8p8p+f7wK0WZoz0QvOMtsa1ZcBV
/qUSZoNPjCWOLgcurdI9p8q3tpa4noEsb0Z5mqJoUxvGA6RsHrQp6QmnMa7cBOma
84fZ57c3zwxZJdF2gbfpml1X4M+6e5zwQTs6k6YW3Wfnq9IyWsmH+O23Big6uEch
HUGTyn9aZgr+Fdsb6fBK0I7FVBr3k3VvA/hKzh7p0O031191Tti+DVE/W5RMFECS
7U8fDU/KWAK4waz4au2Tp5UeQJ6oJptn55zkB0gMLDWzroTMZcUIwnnaijfIUgsb
sjzsvDHua8T0Vnr7AB907VStV28lYO4AE+W6UniEa8M6gtVT5D4IbPqQqa8o8ezu
EV8FNGLfoxeV4A8NUGMg+u+xEl1JvJOdlhk8dGaHBbEdivPxA3Pj/Rg/2xbtoaLY
jc2hJCduTkpAlcuukM57wMAsRrzLrglhNvHAYkxRpe2T/l0gYPXLqEvq++y+cvTy
yGR8lD0ODLDmptH23EagEKAfivc/fx6zLKCk1aPddcPzWzKtNw+cmS2ZOkflMu2m
wRF7G8M9eysy0JphcXeqNhEbjvhnbslrphVZ9RjkfyK+UPDFvGW+yc34w4MOvTxv
aJXtgQ8gPVEWXFfUA7vk8/usc8l3EYWW8wBy1XnNInqCZlQKLf60ZTH9vBnqvJur
G0DfM1nHWm84+Og6HPOFtczfovm/f3lfRRf4vwVXfZzGCZcGKtPVfqkyQKTTa211
OnlJDaGTIfSM7dY3ugMzz1s3a3zLjaUSf5YrS2UkK9a3seOoC80lAhuAIk+PaMtR
xsDFNtkCRFlF/kCdLRYEEL9f5h1v6f5DJkPF33rJRzNbGHzTBZW44EVDMBZYX0uY
qOrpbYq+1hWaNYlY5pMZ/hDX8mUIr18fUk3/Cukg8aaWvdNhrZvh4gQbZN8X1E9H
vBo3tXKLH/VmJhB4RnA7sxRWXWHtdCTLzdCGZE5oiKMejd1g9CSmhvIlk9AUuQj1
UxdGwpVgp2apLPRmFG/nBG/OfqgxjEJTYf+Y4kwxJBu5tGuuOVCaKfuIp9YbnycP
fm2MMocQ0HfAT0XWBwkemevDTJMvujERQiq5PuyEg37N+TjF4CYZ7vHd1iA+D2gm
1PK6xmM7AR0+x0HHyQVptYXuEkzXfsYYfRgJUXreVm77tGLWAsb1hVjunA2ngt3b
edvr/jGhV+XloQzJMAnI/wRKh62YkLUqjWYItybWqlCcOvNXUFHAnRXkLBqaj3z0
ckPSv9aKU+r1h9Om6Q5BufBk9JFHwo2MXmPCgMwAK3z8dVEjzB9Dv8plC17uJMY0
XVRkLb/VRx5beUsdHOXcvwai94Q4NuVLZQTpsNc0wXn2a+HnuoNHvtI5UBZa91hH
MIFSR4zMFiIuFVN5s3ZvfYPrJEoP4c2YnUc9C2nyziQeXBNDD6vqLbbR76fgBJf/
7jaVpA9O/aXtPD2ZiEm/2vPeIm33nsOs6dW+RkWkXJXVy4gJLfQp6flv59h7qwIZ
1yCeGs3SMOdZT0DkBNEKAYgmdkYew9jajHB/t9Wigvu7dAyiX1IPYTc5/v77/262
NaXsm9kaJnYhP1eC6LhDWkMpGZm8Cwff5xv9bTFL/EzSAdN7zTkeUbideHgyQTvi
7/nrouzKnfHfarms/DzWjNr6cW6gnXI66ibefY+pggDfKk8INuVNKIqMcnDzI/Oe
QbOyPuuz6C6yZWXVVm0ESSAkiQsHnnX8XlYc2zfs1zU=
`protect END_PROTECTED
