`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXQspUJ+S4cTkFjvvLhoaaAADDOuvOKfQ5P+Z0d6NBh+KCA0BxUPKhAM0xGExDv4
zPh1tWgkb93kxmlQhiJ8sB4xOVVr92KdRANeAlFXwKS//c5SwqCBw/fvVg0/t2xQ
b711Wtl9w58RGbQWJioUf8c2ltKKJXqFRLhfQxZ6kYZ4SVClDqR0K3dNKp+R7D1J
cd2ketB8Fw+J+LHve++y7veUoM+/TgH5Y7cejO2NrHFmfFakbTqfmDb2a9VHpy/i
o8fAoB5fK6KsjKNLMAarytDz+eYG4wb2l++FBX4DjyOwiid2b+9csF2Cl86Jv1gT
EhtfFLwSBiGxXENUdZhBM/TjuJraYEHjym0ByNFg/0xodfmxcTFk/2j0yr4XdN+A
G32ImzGH8tUFtP15op8B5jgXXn7EZLo+fU5IQiTxQrtEF7hY0cuBcTjhQRJZInY0
fK/MwYrVo5eVc52XK0pkpDgC1thees2L5PUKFEPIM7wnVTeTaOirZ9TLtrsguOWS
PnlUOpR8Ath8x+3mcZ2UGoUJnm/RYma5ADdwB3XOsES9gU2XSQQ7Y7M8C669P/WT
8gGowi+UaDpSxMpu1Rn/brnQvQ6nC/9mFNhzLJSyCgyYDol0MVZjlP2uJyiXo3LP
wLZhjRREEb4g5keMcNDTY7XXBvSIYCFu3WTGURKjAYk+OaMYNEkX1Y3/dZoHyzMS
yPD/v+dBFacYJBOkxBcpB93at7JYuRQ38Zk/uAVVPEXUdmyN+o6U9G8K3D5LYxlV
XOh7+LxiFiTVnKp0Y8/WIETXz6xkXL0562t17NVUGppfp373YCLqD8Jbts100oYz
zqheRmKjYgx9x2vAv6Zad2xrpwgU3+VW9dQZScRjYEpJ9p5bmBoFLJorBnBTGZSc
0icieK+b/3dN2NM6g5EoeXeiZv1KFwtyAH9Oxq6hmZgPMM6/sQtiHOHYN0kda9tV
oivCswfB70pddZ+HkFHCELmJbSzRTczIF9jaYNlL/hI58UVD3BllzMpzSECgXvXq
J6eMBs+BUDIaoS6MZKBLWESJKC9WQMLySuNEPSan0//f/lDOVBPInDpt8yzKYWNF
vqQe6xxJfUmWrcZbp1q8jQIme6dM20BkbbyAFL9yU80rJMXsmNaOGy/ftwfWB6Nf
rPyfzucpoeum4QHX6pLa4fmamgvav4rvu5KeApkjs3AhhbMHydu5jVUKqO0tZ3kI
fyAKpultBWApEwQZ/XsA+dG7V33lSK8P5nGdOIqoCHY/29IMKUiom7TLUMEIW91c
wjnMpTk0uXsrGn9/t0/Ue8egZW5GkZcgQdtHPrxAk9bMrXE967NbQXN+AY1Vx1ZH
v1Ni49vIqK+HQM5FJCpU22e0ZDLV8J1SrV+YnQYZJJhH5dRAshnAnkGcvSj/NYcO
434z7GP+TM0OP/9tQxuIHSuy15i8Te4gCB3FW0GUkGDHJtabIRVYg0A3Qe9mYSU3
QKjW1rRC3vdQRp8xbPHSi2J4bX33NcbgH6MFQBq2AkONr83h52THSlOSpp0yOsbQ
j4+LeDFVkPXzcPAv6sr4WE+Z+cnlH2MrP4aA/fn7HOZt0uzJXQrYy1DCidS+zykX
AA3evmBxj+s/u8hSuGE+A3eb/80KhGcLWBtmD0o1DPALUnl7cShF5OB9z/zwGWGY
Zucz98C/SnZxy/CztYkmy9jdEq16jL0wHJQUUIz0yUFl6edb2sCvQ+2epWW04QN5
oN4uq90ReFom98HnEK+nitVrvrWjCrF6ztlZe8RnjfYYsIBVu28BjylO7UdVX0AD
qGJFOW3k8jV4ZxAeN1tIs3Tx3HJ7IHxQYiprApAl7wSrW7uYzfLMIBPOQ5/73w7b
SuKsPZoSLrfhqdkxtPO6uv8rqcysPsGQhvBRVHyrhoH8lI7T+A/XXt0TKn2/V9/7
8FbR9d4Se41D/vyoLj5b2tg64h+C+1drLNhyecJ5ae3aCgDh4UiP1970030tW7+f
KdIc3ueRSJ6Fu3wYrewHBQ==
`protect END_PROTECTED
