`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MVV3ctNXvfm2qEh3uwSpCEv1ILgJskyxFhXNxjMR0rgcRLSdp5vnVKT8RXJBhOpE
Q/IpIs9P9CS7v0R43drU+C+8av5cOzxmJWkeLscP9sKpiUqiVPjx18JrnR5VkYg0
bC8Lgcmu/Pe//CNYcxdLMn2vMWOAOyzQYSoeu6V6KX/CuaEpuA54BgU4p9EEQWFu
b+t6+Mw3t0v5ZvEX+RLfK28q6uzfQKcHj3vpP8Lld9cJw8PdnjYT+Ggp015Rzru5
XuTEEO74S3RpgkVfLYsyFP6IR94UiZrVtarLyYG7Ikb/gmlmLq0rcT2oWoAAmfuZ
riqorDNMhPpyTo4bbzC86GEMZaMye0tnT8UY4UU0FAZ7RJiWY1zO1sii9lOO4d+Z
dHtdzzXvBmXftfJHEawqOIb+34En9Z47J93lTHZrKDpYODV4jc44wpl1R+c6iazh
DorAYj7M/+GvgEnxsGtJaVcPiqPwN4nLyLmktdas37B5zxCJ/cE0gaMPdz24hlaA
ihOq/r8spOYDJSuGitJpRZDew1/YDxJjna/yfCvtiKoDP7Rn+Y0m8BE7pNiscaf6
dadBnntRvaYjVGw9DaiKTzPJ2eqxrDd9/VXoQQ27//dnGImyk10pXbX5c5qIrCct
8gK9y4j/CxADXUdmMj0Zy3B4Q6Jtc22i9MSzwCm9V5j5ebn+cqlk/HAhf9/Az2Pp
Uv4AWGiqj07sfxQPfKzFdhrqPYz9AJDkONuBitZJeLJjhw5tHQgI1oV9xx6k5myz
K7c4Cpo5PoDBuvvjrxEP0KiOtNbicb6kMUANCfu03wHp9rX4fEaUq4giksH49K8N
/vJej34E+L2VB6D2pap55i7B2jqjRvF4Gxh6exfiBp0ngNCIx9wzGTy95vs5lfaL
z8Vsh6HClb4UfXrH9zPhCn38QSUH6EOVYpo+lZQghw5SQtpKuA986bgTR/z/i6Ka
unlRVJzHF/J/w+0h4sRt4CtGwYQGAfj4VyCoqMF30xJ2td17TSqWSX/TLK6X54qG
8W7GBXc9TKWh11lPeCAujSk7bemn/uHJmU6mGwtPaaOA/OCun1+9r7mlQ8PST8nx
VfRyB5+JbmVp5eNkrd5alxnhzJ5khrt177jbrWZcTxCc7an/PYgQxTewARq/N1dQ
PCFbivBL0D4vas+gD/qxaX8zPYs7WGOAiZqp9NFBlLtZelVpkJcyFdhwBQOlAe2k
/aw2yleoEzhFHXgbioW03Zuf9J3hZxnnlHQsePO0Xg/ZTAIhoRcmtmc/L3QTMeRK
7CRyY1nM3IayWDBDyo3rxn8B28SXkqviIEMrI9hVkin5KPAdO6CK4NaOEYuq2LFJ
hiWkV/Dly2S3exEPsAiih75wRHMhNai456eLROS4tSnsnmbC456VBmODWPHXPl0A
lsrvsMz12dmpeChRFAyNPzr3Br9/qbkPDHMUZ4QUyPr9cthBIJBp0p0i9suMv0qg
fg90xDiszXItA1Ge/4j27v90omQqvjYms8qNgxkRzUt6lyuogOpNr4UYF3g/gU28
nfYePO0GCLG2nDbvDXooxwund9MKiHWR+xO9G2m6E4/0Cd29T+iQiHykknVLTenw
jkHsVzQdjsuetL2UXd3EoB1oXC5L+kRvMKP8ehFt27Kmkeesl5FPRID6Tr5GmMmh
KiXoNraCfZ60qI1LOPyvowhZ29lK+w/TlQVQnoRF6U0i3Kq99iINVvkDI5JwZYSt
J41cPNqA0Xb6Ysi9KoC+e+uUsbFBsXrcsONh1mQy1PYmxkKokdKoyZpmWurNXZS5
MPZHo0IFm7hejW6PDpv59wlTvMi8qv/tQ1AZzUjQBip0LLVzfSJXTxDY8BDZsgUJ
RVYVRci0JScs/AnuTDYFSIjzCA5oDO9mNQvqLp1xG9ZiUFIS/tEKNgEyktj+a21s
B/3QW6a6HH3YnWGcjy8bqtWbZtKYdhvD3j/BIIDLp4PFAb4IObbJFGewqvVnuQ/k
/E9QV7extK9mrtQN9HnhyFVaBeSv8t+/X59ypz2AmH/YbnIxHRVOHhXFnudY54jz
RbohOiBk4BikfzMwlsks0c7MLq2NHaTmzomGX/iW0kfdygR/Pgg3Y5QdsLYIkZwv
Eikr22hUbH41htlAAY0tboBc6LAMmzhyn97ln1C3B1N90Lz04mf8AYI3G8Ts36J4
VaZJCIvabu97cWhmp9US9qk3ceqKay0hQSDp4Yq0IJkI1vhPhkSgKLSmmSzf+pqM
T4aFgSaDbNqoJfnWj8yrEIO9ns706O2VjVYePSRI2cpi0WPXfQNbSP4FTA3h/0bC
t4gulfq9tb1oSoGfpRCzFdqwJwpElglKilOhAgyTqsNZGodoSjiqkxy9n+jzV5ja
X9qWAWnNjIWAM+gRWR7X+BUHG3ms9UHISJMt1Sg81O8Fq48/ZGxLu6r9cXRDBLA1
Gtps3Al/mdEGQAlPsKEtFTtWcuOBlOUwzKjEOfwSEPx14Xt1xc1nV9c8PGyBc/fV
YMvW6SRScWBmEK7lybY07z26pT0PJd9rGt9GXb9qs4AYpO0uExjvvtu3/EJSVJb7
FpXf9N5BxOfElIAus9Ohgg2jC1r3Vv+tZ/dMRZkH2FS+ZcRY8KqEY1rOsFAYHo09
eyi1PzEMK19mn5jrSdfAzwQ5zbMXYM6rYSGhwP8GVaazgtNhNTRi+1RRs+ulA6m0
2lj6H0A2/kBmvn0q6WjlPc5YvlH3CYegWhGox6TAbFtydC/hxQwrdr8hgrSdqk4t
Y9DLVC0fELz/oEiyJFzkgWGSTbcJCOi6Od8cEpL1YnOMkDYTrs+bUSlPyQ/5+oiD
8pew29+QuVSMy1nErUXYDjTBc0o27iWVXxZtdQNzr6vlICW212yZYPWE9BVbOt1V
jg1yHbKMzC2ium/8KnD8y4/bOpKOWYjy71o6q/KF4YDKu0xN/YlPH7BCj2j8xEmj
oiPtq98m2OVZKbGEcb8p7CPzHBZDoTSgq3psW3N+O16niP5EADytCzw8NzZkkiF6
pQQtUe8eBgbPQIBC39qaEoe4H8UDgpdShXUPfdJOJis/c6myavE4PkggnKqMg9Q7
t3p7A46pbxDqlWPe+dc1mZO87Tca9IGtwSkopKeyltBUIsul+bSKSbyskg/I9vnM
NjLZATwmZ3c42f1hHWfbLXm2dw5Thrw1bH37QQ//0rbsFChb1uPtAJwF7DaCRo5S
tn6ykdH1YS0MVV1M3HtfmE4ZlVvq+wxqPkx1aN6aRkBY+ljV9/J2qN++7hsdLFhD
zgOFgrICCQg0yt17qROKbiCS/qH68g2AJw1lYY69zWvMQCsHUgXvJWymy/fDahJg
taViriiZl3VXEZIn47vU8RNZsw81y7F6LLLW0tZdhN5dYExMC5nmkidvgr9SVyOD
yNaFoViknlOhKKnL1wer7sAAAZouGFlErZmAlS1DeJE+JbJUf3VDHUU+GI0rz6OL
u/3IcGAh/YR63Bp2Cn3EkgPjhGvCnjlGn+ofSAOIBfvw9ak97bUGRR1cuWi7Fahc
iahj+OWgeaO3KG5MxSZtZtTjlVzUiGkENIwMFHmN7Zwclg11S3HxcbI+vc76vjn/
I20xFUgD5tNIlQ/xQ6XPr29xGiOBB67tQFsiUrUx/lAhDJ04hmYLlQi6xTwD0HPI
XKznWIy8AY8wnAUy3t0n6rwOwn8187prrL1QhS+S6WsGfNXfHCG0HLoR8I6vHx2g
0wSqlPVeMYHhUQGjDhg4Fi0Rgi1DAdZh2N1Kp4Db7XmAzcCq0Hk+7UnZIY6QOkmZ
c2VAm1WC7HPmpo5L7vDJTdq87PXq+TOZPE+ONNiY5IUAakHZ9mAptTQ6CnMh8f0z
cqs7mhGGLJ+cnvdGj5Enedj2gjdsDIA2zAZVKaKAlrKRDzxlxlrvZzvKdEdbMVIf
uGa1w/NHq78TbNUs2GaWPGh0+LRbCCSRvgPPc7IPNnEY1vnnFds0DYDDJirjhBbS
caBb8TzteKz1OGiZuFU7G+l/a2ODfIQeGHD5i4Iw7SEcW57a5P50MXtQhNjB9TCz
h0hDZLfhpUlMSQspuaPXtfNUSjvHymlK2Q3Lq5V7Ue7YgT5UvUEwXJWR2NXKvm9K
C3yx5E2vSyxoTM+16XAH9IFC4WiDLqZGeYWbMhCG2cNw8BpYctKKJPKKbm7GddP6
+Zw8uarcuTYVzzs+0liCbVJzP0vb8Bd83GKyi2aqm8sd4m142OvIQDkqiwXv3wJk
bIkQW5JxlpuWf+IoJLtChRxse9Gcg0ZEsEBseT5dJo2kev3iVBM1ah+EBo++NhTH
W0jGFYBo7Yv4/d9ymhjrAvBy2gvh+0skLFhzvNOUM86PAhkdIdkrrt586RooYbCd
U3OzaaPMPYABnO3txcrQX7MaXyus+MQ1yzHFkDoi7UDEm6LZMl0ywytLyccAuAaJ
Y/c1MIIV5K/8OIcUugxRGYagZGpoHOdribs1evfks/eeTOY72FGuYCUVVUUkQKsm
0au3sSTPdiFYY3Je6NI2MTwjC+UMvBEk1UWv08x4TtnTvKb2IZF2WVlyMuWK9FjZ
9I4VcA5MHd7VniTyk7T2KNs2qvJR/Ka4eqCTzWJ62IK6jTkS3NqwupfSVfMDvR8n
ExrjLDyTtYzXHBv2jYRG2qbCS63CdHdJAENWMnKTSTNaTZEomi2135PS4c8N191o
Zm9dOkVOdT/tiR2PZW97JATWk9sfntWz4mFyWecbG04Brr64Wogt4dKPzfEl6Ho4
7v+jepcCpLHuBTy158ZLM3f0uWTLomHMQ8nJJ849f5AfC/Ru5FsVjHZ6y6ZM6MuR
Hru5eHErluz/jbsER+5BLwdwLu84Li9y4gfw0ADim703z0Sw6pg9vgvRIVCDbZ2O
BD99VJ5GG41AEashse1556VuIMDXUi1IOWmQHSm0XIHTMZpEM8qhpnF2WBaj0kjf
WIm3sWgV7JnpeahLvNAQR5koT6v2w8hfjvEdMM9fEDFQJZ69zdu/V7D5hV6w7Wz6
+BHRZaNpg5Xq+7JTqV5FO6odpiNzCRuyZGW/Rz/I13qh8+7X4QUDmIAE1/FaXs0Y
EWww6PnB2rRM7kJo3g+ByVC+1A1I4cDi8ww5RLBf8yG847pWpC4uWHI0Pd/gTiWh
gJ+zYqiR9lcbZQXv0VN620Zlg7fxXlLkR38SRSKhluK547zOgKWN+Gy3jVbsw+84
3d0zH/f2LuMCrMRHWDSuC8yA0fLGMrYM4HEKVa4MlsGsAy3Ot8tiDEUXVqGDn+5t
U3pnTmwDb97bcrLmqNW38YDRbWanIggOcZvayIq6iJStq+UtYX68kjZn19MIZDBU
OxpT6i5rCnIByl++zgUgGBFjyQDhzdId0hv1Qv1Yezu8lRB9b3t9wVROYKZILYAq
+jasrdxX40tM+aCoddmQXgQn+0DeMK6GpuRqHssfuBTQjeWNuYYcTgtCO/NTHXhm
6U1bn0VLWtrVzt9dZCsAN5r/VZgQilDVXKwlX2EFqgiE1BtEiq5k44WQotomnRzN
oZ3IMF9bfXhI5AECsGG3r4Un41WHuRwwV6sM/e94vx9H5XQTqO84R4Tif+y3fw16
WIsCOnEnuPfOkNOn/LheZngGNs6M9YtO/MyXkpwZHcc4ksu0YbEtFTPY0FmMQHYT
e/plbUCMzrl20jdK9h133wksTFIxj67WFmUtGcdhNCYImbrYootdtKaQXxgxKNfE
P9575JZY/Mpfi1fvAC+BZTbGHBl2XN5jPSSmfHUd59PYvZsy2azy7sus4kOdW1QX
MH29imYjrsww+tSv2XPtUrGjjKSFkuXnu75vu+FXno+NNITjO6nCrkps4Mfxzvvu
sz2i5tFovemjFB6BzmPeAulxJYm+5qP8PXjLvoyQoxzNhtyXCE0l+lgk70ci3t3J
uXjtbdLENx3CXbieeBjLoZyDay9fQoZ7F87zwM64LdTvhO1YXPJN3K4sAaWuEpKA
5So3VmrlfIvI53CPwoyrEROR0cWT5X1k8vviWalDrrjJgqWl+tyST88QKAnyM9M7
efSkLfAXCH2fhLqfpfu98fP6UxrUHR5mHCRmPLZ+jaM+cFcedFKVm0DXSvfeDg5K
XcMkPj0xn2Uvbp0rGrXMWMT+dyXLUbuXDuAO6gdLtlsDn+2PkFHf5Bs4nsNjhh/y
+vAVfFq6tCHy1isZBA6fxPRR9KIorB9xJ8TI1UAQj5Ge1C+hOlsvwJIuo6viR7wX
7sJCGWeYYZnrnTjIThXmLpBN/mH5PV16reQ6/dyYD0Tq1i5z8RxCth8OLRefrXlw
rPv53b4tqzf0/j10OxrX+Ybla4tUxetpZWS3rQvxab6br8nvA4dW9CA6Neo64WRM
WWWeY/Rscc1StI5a1lRMsVhSTBuPH60XVRW7oChRnXu/HQIP+7KvooOJgx/AP1gH
yvHPfzy13AHvrAg7h77MJL+AVkRoPYqLJtXLENVrizvgz7VFMBi4z57ZrAmplun2
kCPpY2nE2LHJelm9zlfcHq740wzs7r3QYUB08VOsaUI/JhZgJNdw5GRc6S7nidxU
2+FyG2VeC7b72uihoWQOoU/rCc7nKJLpXc1Vzsn99c9VNwzl9kt9jPTnm3S9pRLE
iJSKDwgCb8NgvIYfilA4Y6Lh2XAd/uarcRExyfFOOf6jPKJjUbkaSVL/qWEvPx3z
tTK77AXlrqBel3J9SVH4SrYZDEWGuzyI4Mixo+oWjDc=
`protect END_PROTECTED
