`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mNwSuPbZmWqOm/E9G2mEZRwOtd1o3kU4tHwMT5j8elGHeyW2S8uei62Rm3ue3ML
5B38aG+Lo7EVFs8n1Fk2zVkmOxldwS5rPVRBi0s1/GYOwLFTRzb9D8tS00p2mLnK
F9SktOae2ZGh4tCCZu/1JHlr6aJ9gr+5Dec9wlWEF0r2T55A2/p5lTHkN9BWEKLS
qJq69DJnj3lA+A+XMDSZck50TYMtS1ja0IWkpwFsDI8wdhwbHIqNAuS4a+JVtz/m
sz2j97T96h9LZUFx5eFLNxdcOTALEqur9d5djzDQ/twhOVBWZm8wYP8dIG6bboTq
oxxgvf2quh0fXjUPGHkS/lgNHTuxexI4+ImbXW+eGaqi5W0fU6UPw9gIA/Qju3fQ
L+SyLE2+/kaFYIqJbhiyH7Q86lcFpzHod1ewllhKJO0HNUtmZEtNrLM3zZHF78An
A+stu6LM++lzhm6eYUdc9a/UJzZD9rnHC39XDkuX7znTq5+G3YWa6J2/kjYbfiye
L4Oh/bIFE5CyhdjZaZ+/xGlzcR/nrfkbd0020muk6JZgMkjpIDeaLj4H6/YiE2JW
xy1bo6rQdErIv01pwAqz+yMfxrlP1sdHHwjh2pCYCf6HAwYPiuboDIRXsipqrT11
aQoGzBsMqFUQbr0XunbjUZYKTGTz2Ko0vGkEQ8joyAHXEDvNlUo+xY0xywycXikz
T6356H2JA6CPMbS41nkGHDeK7rVGL9xwXxPUybsukM/1jqLqKASbDOkWgBQfcr5J
dnM3EE3c8iFdUnPXb5NhekHseorVQtfF9mNEOJoBZA7WtcSRpBqeaMDjnYJ7B7Ua
/LYY9af9Duh9MBcMpHL00FbwPOkUA0NMnNb7/RQRFpz38mDXokrdGoswkWSfPbLa
3QGSLIVquPgPX3WxZKJwJcyCldNB7Ii+UHyx1pbGTCX8CMmFQbXJrxHAN+yfE11X
mrGDxG4n3ewIq4gsk5f9Bf0fqmUTP5i9bWNNNFMzK5Oe7yiY7q2FT/K7DWlbiyBF
7oJfPneUQDc5f/FDouNUK8129t+hYu3yWoDQp7JaCDZF7WZtYgK/S0PSNS3EhPDx
1ngCmYfAJw28gcy5PBNX8Cysc7sTkTfWoMdBerFj5oqXLUbL8PE8sCVLndJgneeS
9OFuoyMeWQT1wG+ZMsKEHW7Iz8OmI04XFyazoI7Bp+tiAWFBTImwHqvVDWHXMm4x
quPH675kIWrR7m31RWqbsz0+vFnqZy/4bUishnX1MQV6HKuUta55ph98W1vZGCKo
z06x40YQ0RpZKhOXcowIXJjeVMt2UY7BAzUkrX4Jbt9Xpw0ERo7UiCpP+a1ABHR5
zCq+S8BA3P9DixcxtZ+g9mHGMnrMcQynOjK2nKyylDW1baXoC6NCakqNFIHEytn5
IfNYkp+G6TdZ4KCtMwoZ2CLIqhnvvdHF19y4MpcEcthAXpY4WUEepcBfWqxehUzK
nYgliyJpEeL0gRfUSg6MB4xhtEOjGEfTDuNt53DcYKwD84QIX/UyqYaKbdYRzdS9
mLd324nvNJAQARa8lcXHZBE/Q8j85NlktuvnPhTf95NPcdAgR5v9yy/7bl/r04kd
RFb1NSOgonks44/opGZ7GGw7OILsz9YZnVqUkI7FgvY0m7tiumyR0Kwz9QroqZ1S
JMSVSMq6EOMU1bogn7WVYZrUsJFS5hedh8vX9kmHBCYfw/3auUFlB+lTwTaOdKSU
X+hXsb2CHa5FhLn8TFIg3G2D8mLCGdwB1E/bW0NfN2RM+kDqX3y3jh8XfUqkyOsR
FoYw/EplkEdJgDqS8K2ZSyc69ca7pogwpFwxu83Xb8m3RkGyiiipuzPXT43n1ytW
Yo5MBrrHmybj3BKNGt8rqQdyXyCqEnD/PRY6xm4iJJ3CIhkxRwuwzzaXzgn2ossZ
VSiyBBsbI9NF1Qdx5PlAg1uE28V8ihDnLGppCWhnxlRyNe53uOQwZeB2EKFQTfoa
Yah4+HY2yn6OzfKCPXh7NYs6Qmh61imYyaNG6EaEy8hTeFjpfNaZbPr8m8du/MtB
nkeo1/4ZpPsIyNl+85CUY13YcSsIWn/xkBFDA/lVAi+nWfSp63Nrlg47C+t2cWZu
q8O7CCJz7Nv2Wmo8fToO5lAxzm2DDSQiY4BvmIhSw3A7Oqdi+KD8+Iq6jot0CGNi
DMkT4svy8BuaAE3Eh8GK690yhSHmFdBGOiFS48YoDqmPswyAKXnyrcHJAchqzO38
+LaS2HRUC+Iqff6bsVlRZjv683ifX24booVZvDFF536rufIuvlI2jIdWRMDOG16r
sk52KKOhO0Ir8L5eqz/A2dLgpj9RhT/TbiIkiFEztR4v0TrjRqrp8l3oyVHME+AY
AL61bHadrWdvZS5okVLcvIEOJ7qVeSqedTvniw8UgOX5OxaBwnnmVCMufsTukBiD
il7hNLHva2wftKN0BI1nlaRDNtSWvw3XW+xJ8gw/M5zXiJ1tqS7lwnCgC29FZRoK
C0rMPpKuotV+Z7oDXkez7/MuWjP3ci2ltMF0cmydtUCl4RxGXbqoK6zoQtqDviRg
Gy73pRgrQKiofj0aofSYwXZYXvn+zr05ny/coBmC8+wxt0seWorzNQryFoNCk4PH
pW0RrTOZBzuDq3pEsCLYarKO6BFxJJd5W5xlKLo83Suy5/atDNx3MOur4NMchlr0
lXItrVAOuFv3QdF6giuDWot9QjVzqS1vUN8QXlGrO1UVg/WSa9VyY/qJtt66jwHp
60o/DYlyV4Xf3IncXHCvSLKtFslKaJdFVR/j6bXDIJSDN1CjyFSXPrKIW2I5jmZR
GWxA+Ww4NKeroHh/UCjTbSQwFwgx9EY+gXECtymWcVzicnpCqOd48pdkDMBpjJfe
txrRo8vjtcewdrvmwXfEoxJx81MNmQ7dTd4kUq9pQsOFlqGYnY9Zwp+A5KSVqt3t
oSSsH+dTPHIlqlZeppYw2mjKLNe9Bhg+/yHWwzotT+mVy67872qIwebpBgM449a3
1ZSA+2YFm4d/l4Ymb4mKvB9mp2rnOY0RGa38sBm1XGNzO8jizjQtYgFLtfG5oJbe
GQGzgDou5JT7bKgJs0/QUkXIhbCMMscaayEagl69RLtf+U3KrM2RSHxpByg1Y689
qvC6s4OWmv7mI2hOArvkEg3jR9oWDxblWmAWEFOh3GQIPyTM2sMrGFBIq3TgDzII
ISnphinxyQWc/I0oG+7ZU4GiJ36IvtsvcIKaRfjiQsPbVM+FKjuGtYNAdumb1y6L
30ECFWB5OzctV0CREHLF922AJnSRa+x8yOP9SBl9wIdgdMo8mGOUdQ6xy0PV3uVw
R0mFymj/0rT3ny1CnyzmgeqN9MZaaovDe2tu6WvBlMroy1EPzRNirHl4ypApjW4p
8LjI6MxkBMqhS/Tj86LMFRPigIwgNBiYx4ph1DvL5WNPxlXTwpMz0sIcTU70Se2C
9XnmDp9flivrBlv3XL9f8G1iz8QFWi/Z5cwHCqqrjazi5NlXjy79A5cjyrRE0nge
1HkYQ1JTaD9vQysAny3922fVF17ep4jaB87Bi6x4mWQA/aVQt+Pz20KDyQ5EE01G
RLcgA6s/uTILAeyQiN/43CHiBqq5UkGraldgXZIvKkTCiaY/XT5diX/3Z6hQQ8u7
5rdxVpDyLDbcpdMdQ1x4WElj7A7UCeGemUcL8F4sBOLDcGv3UP3nG1sxxe/Mrm+T
17ShW+jjp/F/uZFHylMeIPYnIEc+7nKhwM9uoCTT2s7ghih53E/QI51eMfxiXE9b
csANC58mZorIWaNSXwCGYkM6EQuxaCANpsiWngNm24WBK2Rw6XL8xGJSeJSTJF5W
ijMBJmGtrY5Ej2LBGQuvaH0ZJYSrN4wZqlGcTK1E4xDVax03rlQokeDb98QFG062
/0aRmA3b0ZUR84q/nPUSP5aIUWZ93fDjMUmNeRHQ7iFo4E1hZ7P4oqQghggdWdgi
+3mZWg8QTZU7iE/mPTAmMxiKIvpgr8d+H27KXmDVFbJtDybxV88qM4BzkIYetpb1
5PGuHMyq68Oacq5dY7as7au2B8WQHaIULLdXPAU3kCNYYksnUBkEIJhAjoi2u8UV
Z8gC3TDhVlhnxHZ2XPNGp+QrsV1N2YCeZUjqCqurGgJ4UMR9G/JUm4Ww1QCX1arL
TarBwvGs3wkrv0EKzKIIvSBnbUQvzyjLGzPzUwKmHQ6nypQ/qnQ/6dwCXqKoRinb
6b97sThWiAfkRoFenSIUV9LthzXQn/+U4fDLeP+bcuSeslGTawwMvBsrvL1dJodx
ZDc29Lne4tHVtkHcPLLsq/lAUp2WAvElk9TA23TdNBUosc6FPWeBf+pCafwcAF0x
efJgw7EYmlH61uODtOXdWkCgnQ4wzwSdbAJVTh4hb2TPB6d2+Y79Fdh46CbbOdwA
hRey46kFSBltz0CwqpV8j/3fdn/zRByLMLVP+reOCdV7uIMEdc33LdD/0J4tXW89
B2NrmMZNgQr+PjkDiL++BKNELemg1GSPgdWlUU0zSkhAZlUiNe4v5gDjUClR7BSR
zjQmNsXpWQ5sgqIcjRWxIvVkaIZz+m4Fop274pMoeTyqoNYzTjJxKrhrcHEUeXhf
pBL8Wh81l+1T3r4tkrxPM1QJpQDQbdOvkFgeZUxU/a1+eW+cmE4KUJp5UKUyCHV1
6/tYviHTmw6SHA+XHf40SdgWmuVaJUakQXQlvJnowgc37RUze96U7HdCvkFNT27l
q1Fc6MSqCLt7ewsrRN92T85DQ0b8Y0rlquPPfH25RWN8Mqqm1SlMsHljMyDRLOcA
gayISXsZzLMQwYifMcNCnDBEU6YccUgJPJWmUnGkfIugg8H5zYKtByHgOCVleODC
SgqyifaMZHw1oiEaneX/pM0VxNP2KmXpstQulIv4eVj88eJZ+elgEFDCyknJCEEk
Cs0ZgMf+/r6RsjMAYXkSJswveJE9MNoCmJk4ua/GABQmZAjh1tnoj1v7h8muIgkg
knVzXDy48FlSuQF2ZU3h/qanpHPTecbNGdG3+05t4RqFfFSsjwCmCLGp5yQNG/XM
PfiXofPy5l596vSRWu3CViT8WHfQdwwvL59G+qg/cdIktHelukaRjoMGPYKT5WOe
47SjK/XQEW4ikgzwDwXUdR4yC0UQ62+mU4bohrA9r0KZQA4LpPRyCTVBSgdxjAiz
xA6ExZBJGZAyzEWzokIAVTG0qN2qiIVJPPpwJPMsbkjy/CxRGgFIsL3Qg3M4PRCX
BoK5pDHspJ0FS62hDhGSdJ5RJP6Dn6jXEExp1AwIltdgE6J0xUvoT06g8+y4qhz8
Bd8J+nPWcgFfVU8zrP1ynEOYooJGroSo8Y1l1ZfAGE1k3z5zfAfmf4fdBPCtv4CX
7945nwzdyDozuYdJjzvh5il04FUZcBWtuXh9JJhJ55aCeFFK2/ulSo28cItFZxKY
R9Yk9AeWUfPQ8e6MiIytoqQwyOmcLoT2O8q+DGIOFTjekhngvIP7G72BXNGJXS0F
fXN8e69rlA0azyTRPE6s5sfxlta/Yh12bxhJJFy+O+oAUUchwJhIcwX+d14qSrGq
O+zTFNfdCuYrShQV361ZJv552T6uDPqy2bmPNG/FkxsmXqXOsGk1dWCdDrM9M7sx
kYRTWxQtC6Uk5bDlvw1qc0sflBnRpXo+B/AdVr2mcd6FOpmOrFQB4T7Qlwpg0xLM
`protect END_PROTECTED
