`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3pFgXHpQhl28Vl1AOe34Jx0mmnjab94y5bsYJlxPIEwaOxmMsMFQaYK/9JiXTxoF
8o7RX1vnOswvPUPLKHnJpKy2Mmi7BQs5xxV2d0Hq4T5wPResNbPJueIjrtIrfzOh
mgGzyCskOzRSlzH0iIvorOCIcMen48dEO45zbWQPPQzmxtPrbT0XjPfjph6w/gXv
TYcqxV24hjMgvd8MRATxkxNljS4Pcr2SD/kjsf/pnwvzszj7aOG2wSaP4q/pc5d2
9btFhbe6ILNv5MKh34LCDNc4rwf8uBkguraqNh+F37pGPEAVI/q45loBZkihzpxz
VJfmSEFwLELS+HXSKOtkTI4yC+AbgWGwYR23Gp1YxzJrnLyLqJShaMtw3bcd/Syi
/eALIb3BScEopFHjVGhcBh+mj9K1rEIFqbK/wPjwBIyC2KbMFSYgMdyR37VkMSLq
75fSrI22ADkMyVIYsYSA4anjEK2K2snGvfDc7sXs4a43ldw0OBD6V9L/qdu/fYwg
XV66ybtRtAF+Hh1psH6bgUn7kDGRMpVMEDmycAZ0IRaXregPFGeyYbTzQiLwMJSo
tuGA9uXTMeJYLSM02NUvc1WIeM6By9EThfN1AMhBRRWGcBcxBpr8A/Nk7YrEc6Wr
5a1dCxMW7/3Koe9r8QDobLoE3sOCZZstJfQL0z7hOjpjMkNbPGXJuO8vZU7v6DsL
FGBk8FhbERGTw1gZbcMx05id5a1PHd+fLDbrz41N5Hgbr5CKUlPBR16eprURvukR
aBhQXv6pl7KvfOnKpdzhuQ3rS09rmBXNNhfl4b20xFR+V4kOsp/ebFZ2KL0+XWNI
zjEkSjoggbeMXS3PxY4SdC0eLl57OJYuUH/yt7zytQw8Zz44zrbqdOMvpuVp5wqg
tIRccieJpl34VB7W+a0trKSTlkkzAxEK4ZLTHIXzVpYzzijDJaRwQxqyJxbHRsVf
1Uaaet0jVswy2uECbdJEmOTfFWfFwVZe8DbwRNb7GOi3mpse3gfFrjfv1XQEbelK
XVoyc/AH+N9UjCNwUnkrbENEK1p/5xV05WHKZYKFNU+cUL+9lXPQUpZjPg3g2EdA
DkneAcni6VvsoA2gaQQu8v3yImFmuIRdxKgh0433tfefi9i9C3MRA8wsnwEcWbVg
RWry38AmSviHocDSzW50uoWwlbPQ+kYuF9JWLxjUMjmFvmFQj8Cj0S9Vwhif+09r
fakhJVPg7SaIAypBtgJM5/Sf9VmoE8hyz6l2vxEK3ZVVtygd+tAjmIBsj+P67fAe
cidElAqRM/4+EWgB1Yh6XnFQnnnaKOW/doexm/dthobrVcXeSZb+7FcaGXXvjiOR
2TTsznxOzKK3BO6gs74119biE+Lsc9VtqXO6giil392LxfyTJHI2qvnimqk2FS84
z6iVEdkymT8gEnN3sPVNRagIhLplw3605ruMsI0tj86UJYx5UjF5yJLwp+WuwXrJ
8OZ8SDBbsIkolIaZFzUbjAWW9SQSrTDqrXulGtK4pjWd1vwI3L7V1+t/Iy9H7TdK
L+K6EhTK4vXzyP2eOjzgCdQ2tHd7N0z7UcYoHoa6YL8fgikfwHoMNGXK52hypMPh
ZnCdSV7LpJ+xK52sq7xGFIsR7VGyg90noGoo+SUf0tM551Pva99To6VICm5sYCrV
f23o+mft4BXGMaUMoa1ca1EE91JNgBptTj/JFTBXOS/8DAvmqK1H563u4B0WDj7k
1v49UKGL0eGDx1byg7G/Ac1YltVXQM5ZoRWRyztzza/ic0SYOyVWeb55x6Ft9Fcs
mXnEz+xZtMeopifprsZhB3iiQZizqDCe8/yK3tv8p7Npu9oqmkaQkUDDmGkMFOTk
zG2BFGiUKd9XAOhogaQV9JZlyDuSzp7veacYBn9LPcONwurhhuobSU22j0V78lZ4
F488tq63nrcSOwdaMUm7+Z/jlyRJ8zRTvqQa5gzpE/lzv6HzwJUGCR6ZSbcQRFWx
SzJ1r8SZsyRVkd8zQnNH/k/jQnyGA8RUBXcaj4OdT8pEE/liuz+GFZLOW9/m4csx
X6ChO3pUZQMTCkCk2AgYhA==
`protect END_PROTECTED
