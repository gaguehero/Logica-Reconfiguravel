`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+pSeDaB4WdYdD/1v9nrDiOGebNYp2wQDD2WysI+eZInFIdhuUQrRGYHLto7NT78
SmlEviqcNoDCXofeXGNRqV96klgB6EWYuH7ZfXaWX9HFZMPgh2CEarLmu/PwWbfU
9LFcLqiULX6/JuIOH1YjHQVXFgDSJM8HH+ErSflyDGBP5WPUxMQoaGMynPd8oR0w
gLx3P5NHOx5cCjrzmg9otLfqErUg78f0W66daovSvi0qPDeNKa6GQ92rXeVSC09N
BD43h98gAXrL1S9oj36cTm1qNB4/cH0BqJ4kQoFdzE01kOZJZVo1wBgTnr+HbUKB
SplMuGHk/uig7Vsqdo7BciYeKhMM2J/xOBsoDpe/IukzMHVjFqALkQo26F4U1dqI
9AS00Qm7s/ZlR9PQfejm16PPxNDBAuYEyO88yvK6zetJRXPp4DjTvx3GvtuMjfRg
ubVNv8MPW/vztcoTxD5Q2gDbhtQIqPocW3FkQk7FUwoYpAGa/WmkQxJ+stp5pKCk
jwojFDfDLgnKh5a6Zf2X8J48fRChiEM7CT1Pavr8Kbd26aVYlpVzoZC/16L/IXCA
2DrpTHFm8quZ7mQbiZVctpJAZSfvTPDdjoKM5XcogDcUcxvdU2G7xBwze41uqMGm
oJHSUePCgEnL/EldKcsub9xjiwI1haIDMdYIt52SJGAYkvr5CNpdB4hlPKeCSox8
Oz9BiGVltlqwyeD7VPckqHHWKR6PAa2IeswrXmME0S8=
`protect END_PROTECTED
