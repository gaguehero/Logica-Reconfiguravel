`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQsg2htoF16I8gLxU3DP6jnmZP6g3PGbHkegcBHoFecfoghbuu8ujUzhqU0AffrZ
7ypaNrJAgD8ibQsW1qz6PjPjodCflMnXXN+sFk4GUk/0EpBC8QnAmGhPL4WtJhU7
Ove1Jmr7rVN4zcx5DS4wkafV4qNACK5mBQSLK8rXmMSXffZs1yxh0fBlRLA05yzT
9yHDNxZLDSLFlQ08vxqaj/r83jaYgwWCzUnQyEThbWyUwhyHzM2GfkzMF5UfjmdU
iDBzh0rnKNzRKayjA1dYj2g3CanaOQUe4+sAExJX8ZeOHLC5BVxRFtolry+2A1TK
9FX53+4eVL3kBcufy7ckdsJL+GxVrVtVNMS2gumb8Fk89IzMJCgunw96JVdctEmu
u/7qFpfTn0mpYvsnuVI7Gxyk1bX1qfOF0ak4VnQBqmXv+wFhohmToe1ZBnhJdfqG
CgV9eOCoki2hHprXuNiZgDWMoKLgoFl/hs0yBbkwJMiug7mi+E4XHaR/q44RaEoj
ZV4wopxBBMgvuEAFRmSju2jBHdNZ/GlO4kPIyE04pj911umXp7LACW7c0PAxNG0f
IjzH7gF88LXAj0CbEJptsBszqnv4W3gm2nW7zCu/b1zOF07KTtgi3eq4wLEclSjn
0UuwluIT9IsgFcGRamdMuLcW8m7/tTwh8/iaVGs6UH/HvL4WPrrRkpN5/tN9opSD
BqJ4IzAG+YI9PjdCmlOCOiMEArTu4y8Lu10bMR1iP70=
`protect END_PROTECTED
