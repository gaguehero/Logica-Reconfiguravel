`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6o5yEHQcduK3cz9B7m6ZbJ20YqA7onZJZsyeRPDa9ewU+UuD0OXAFRWWnf3yNvBH
MiT1HnWL/3GqabiUE+DVpydMzNDrxnr4N+sxCmfa+GnORB7KHI/Fs3YmG7Q8HUQe
3Iv3OFzUIXGRBL6+dGLN+v6/dGpctPDUhtgI5BLtKkIhEp1Z+21yegw3YRTcePbI
7Dy7QbC/vMOlieJ619QflHNYWyNHeQ0cecpUEeZ/H15sG1hYgyN7A1atDnQNftvD
LRHoSKmb4FZsBFATnoJweeJ2gL1p9GgSnggOVkbXA5wbGsBXp3nft3snrFl7Podk
AHizR+E//FHEcyCCmiM6l3HVzv98T+4EEd5cMKCUkdZsI60I92a6tAKybkDvvq6J
ZkSnwHvwfzJGpp6ZZdPvBYQvmdjYltfvUwAlwEQT9pXn1HSm50AuQ5olpVOEghty
4aFSku7idN8VjGkMNz1PTjMo/aJayCrgUi776+cyLt1sP4+bXHzA/Wqa7y0w6029
WJzbgXkyEPYMxs/Cu3aILyOlheugBeopcX0VapJJOMqFl3BQmxyVrIWbvhQ1s24Z
ksaR2ICm89yqOYI9KV35cIXDDZ8jAnQMH9x/VE69mVD/oYG+gm2FQY0Z3oQ+CVz9
ytA2LL8dXJUz3oc1pGMPTl6nOb9oxqEoqTb9W0Y63hZOoNX5zegj3GhXfMDKudu5
kmEfpnUQcQ0Ok5NV3Tg8PrJ9/bRd/cG9xGyOYk4RjpHceMhpf3/h2B6sLy9/zzHR
Kwj1PVfGoSFdMJZMmKND8Juriif1TfsZQbT2lzKfHUDo52KHT1Z19PXaDj66Rjeq
82iGs6JbW6XnUy0nOmIlibXwkvqmYK6SvFSeHR0qp00+YXzgRQuILtAoa6OfyCmG
J2hBy/5ysmwtK11WvCdEDtpIQNe+d5lhKDulSwNxTiiqI6zbN+UxF0SF1vipdE0V
Mg5y+8sjsZ6uLu6n6KJnVYSQoBfjYGjEjWGD0GO230VL3HkyTlNqI8JuY2GCj3dz
By0FbuxS+mwGPnLAWCsvP3gwrgL4MD38yS2QDxOjd6IjsfoHweADjntkeuu+XFu7
QHDTVP9chUVFA7JHN0xr1djKCGCefhIUrnyGibX8xN2plBaWbsCTSs1qrMNvsOxm
7yGxiHIkMCHaBEUDQyvKxoDUfM+RBF+0QlnlSqxk+IGUMXwXXpFo0T9IZuZsjH66
pYz+bPh/6NqpIggPjIoEbkmHQKKYqzJyIvxsP3ZwjYT3fgOX6fasPiMtLnwrtLSB
fO1tJKdZ4+t/lzVbj4gYq5rplA323YhDeV4tK6m+0fP6RF5zGqlRB88AGKWG6Drr
hCBUfxrfuPD3de2igWwvBF/b4fHKC1dVJaljHQ7JvGGZcsxl0+ZvFOfnJ/9PZ8+g
9c6p4BoXdpqBCpcYm+ts9Lg1jc1MMV9XFFek6u9cTGGjcST1Dgd+iNJc3lhULLQ+
8CrygGpAzk7jtkPBnqP0+Hqc4fdWdyku1KbZnwHaXH787nA9DMhL0VN5mZtJ8QXW
Tku25lOC+E2yb3hFLks35VlhHKSt572vVhQ34zJLMCmuDMlqp81auO2oeooVi//2
a5lh6rAMcOcTdBH6m6khADyfdsxNgKl7a3WCE70VQCbx0g+UaVlcc5KhxET4d8qC
SgR8dFfA+HYtSN0kAUBlY86e0dtUx8ZbrWyIaCMDurnH1LOyCbN7F7i9r8twIn3E
tY+tfto0EMw/I5s0puD4GrRhYYeExgSUgfwtCNstcu7PptafWuTdGP2utkDXmuxj
zzAE0LGwhgyMLppj9qNO6mXOqJF4MDw9uzuEuBwsNZ01IrqxLNt0zttLsm2cKymc
eq7j+tU4upQyxpXVtBjYc/mXLTb8OnRPrprlF70IKa0Kefrr0T8qy2zOYVDQv+lf
u8IKPiLprjlmOJI6+9oeVVdgbWyo4jwHanvqV6/ZKurriPlNryRBNmqVUXFXYwDP
mx4lPJR1+vRupbhQ84nZcMvXIIFlWGXii+xbWyfftjjNoBf8RK5CqKSPPgZgATBr
dwKlDlRIyICcCZDkrXeY6xWTxwyjs923rPOJQKsqk0l8ULiFGO5sPH4YcLPav3jC
J5ek46TDlAkTKv4IpepJv+uoVfe6liY388GrlhnrFHuaOgPnL4bSVNQEBIMAneXb
en3/kehj+npT5ugUkq/JQzat3LtChFJwLNCliaP5o49Rei5eBw2CTjucVHgPetX+
/dSeOKhnopF+hPC2ViBnhqqmiYYNkpHUdOsn0mAFay2w5+UgSIBqWB9rWZtI+pxj
fQvbW5ea6pzK8AofPCi5Vt/XqJbt94/6cX1bEWi8lmKxAinllJk6/HaaJMtMpMrf
1WRrdyMtH7+9ouXDM3k/zz0/MhB9hcx8gfwyFUIdT0hCiOg+ncaRn0dXi7wtNaCA
wg01JLeud6gIvp933VxQQ26frVo3fPxOyEGI/YaCKv7AVBHzHNRcBvyNepO388WD
rV4Vx9wIYulywG6iE7YV+7vFlBhdUyx9iFp7hUHoqc/zspbjVPhWqD7pd4LCw+vi
w/KqzBPonulpQM3+IJwJDUiIn4wU0loidJ1b7Aa/DNpHe+Qe51iQ9DBXg54pnDPq
TAw0al97cp7z1OPEFIViZKvOfpzc2q1KEGwn6gJyA7aTRSdnt+LzFc4Q6+zjgCaI
11/KdnldFpb22Dnl+lnC+hF1im4tEisgSuoiqfboe5K5WRDeUSqFJd1a2d5dZywv
ngWy3VcPf1GriM+5LZpksKqymZFkmiD8AT5RJSMkIMTtmYf6URdHA56hELGN/Yvd
JtLUprRcPSE+ct3+8vEbYUQKRQwDYjT+L7ar/a7GbBiaxcZYmog2eFulZsiC6Tpa
lfDsGcWRbD11/2t5zmCj6dDKJtoY3lznLeRFuyaYvVVLqy48fXnxWy9iu+Am5iuO
09lE3i1Y16kgvgAVGqk6/DUSaJgrdcW9TUAd9KdNZ5IfXCS1sOPRGvXvJDDLZqG+
Wo8ElCnAtrU0cdyKrZ1K6KtUbYGbpOxzMyj3wrfxo6PhILvfJchtuTwMryNiMwkn
Z/sqZ4YPCI9wrzhVlCQxL9xsTD3A6EAZZVsAPD+sWUC5LHKS+w/2p/qWlMlMbUP1
9nyccc/wkeiYOnqKZrobAsLpmk6S3fwgTw1s46ARoNWjlOXSYQk7v7u29G5w8p1m
cCI6XajI7qckLZm8zj8wFv4W8g8J3+bk23GfT1ZND61FhUBUtfw2yoQg6lpXBYWn
iQTvnKsM9bkVsG8FNB44F38N4WU1/4KD7Esw3w/BFU8I7YsgB2I0pZs9ovRdGwIl
XOVrt1ZHTyGQieZqRL7CkXJn3lbUqytOHq+awyC7HKfX2e193zqfRtwQ++yZWRFH
gvMzQ3iBI34BqfA9B4bQE3hQoEQyv13yakdkZ1kgAW7kWX7AsloUS48iMmQ5kTVY
9B6nto9CKNrK8n7CEMGMn7bFfjGv62k921NsFELLloUrl/3AvsL0wZULhR/7JX8V
xHn318pe0nbjBSuW3g9i79jv58b7WnSSK0bW1Mo7N4Ie1mwApzjLKIAXL5q5yb9P
qXmYFDVHJJ4pJLzfUjnLSN/53ClFfz6t31+IgUw70jOexxFik2wttepdzbHqcdPs
OPydwnRXMrtWpwRMbhOUP/XiQPdTjznMIWJze/AuencnP1FS+1JHyMeD8nOrJej/
DcMdLh89k99x3zkkDQ9uZEcvfEUAE+GtXCu7CcaZWuJNakzSFOuppbanA9ssendw
3Yq5xKvRux7Qj36qzacvPK0Pxh55LhlLAzNqdP+gjDQGQhusSTdSmo1ifIk6JqMY
/ExByxExRKRBq0LZnefuq6der8jMfVEOYwi/LhGMimLDfF0GBUWAqtWNQhBk2x5A
vMnj8tqbpaMVbOywwCEJ7J6zNxJQrcTOIlGJNoRr/vS96fMOhCGvosY9MDDMDmpm
kYMrLEOleKSwCsdXZSr+HNgw0EO1LcRakchyrE8tuQZVYyCaTfvC871y76FsDEtB
UpJdVVBn3ht9wWMg2HAvCgf8jbBxhABdXlSiRIJ17AFloPJtWZBz+LWBgpRC45TW
1X+svedBz37HiioD5JOEljbJWZqIHJF1ieMCAclhg2nWLiTNRKyfvwgM9NgJ4DBy
u7xcdxD+Re0jSww7h5EH9EWjXoV3rLeXIBPnNge8Jf9DARclWH3r5HvW46vuXfA3
Z2T6/UQJC8UgLrr3VGA6pPFsyno9elSuFQYfuZ2cDZxG9GRLncnHCFsRmvm2WhYz
AjFrE68x3biU0Vstgqm3Dp/u+VGdIFY90xliiAMD3jTjEy1EsYzJ/7JOUD6yEb/8
WyqrsCMkjPPR9c8sLQax538PkeDGwt58FEky7Iz+aXSXHOMcyNkjo9yHPhDNM9va
XRmf/it3CqDKgLW3PFyjoM1EEGlu0dB69koPBjmkpeiH/Y0KJOZZx7/3TnNKc4Hc
tpbAKiREoIShoe/OGYNCg3R4kakvM85wkHkBBCiy6i9ElCvzoX3NiON5dV9SFbAc
xRntCkEh1o4q0COkuNl46NNGn/b5/CP3NRhMD2OwH6XyP/9lOLhBxbyx7H8dI/5y
mexQ0vncNrN3Mnor8cB/iwRtmNA5dYD9fYHxmcvCON0lY+HuwMEY79G33QCuVJ8f
XAXjfcA9fcXYBEEJHbOYdHntvNLL/Tm1DzKDvC0pyCtPUvN6AMUw36xjOB2qNFty
vDsuLxzgLgp3j5UKFsLC8VzEShg/in+oUrBdhvK2gUjprIye2818m6W4SoffmiH/
4NHX4R5oe5KIbckZIQVKvM0M7zUVRJq3YZHo0TiE1O3ZQ/Moafmg0XQREiODqRHt
dSBCv1Ejoz0PoM/+lozzKnaKkTE0nTM0LBdd/TAdsV4cPFFe+PqaW6YYNhXEiiHo
4nh8cSlMN+wswgvyG9UDzmLYHeVfRv35IUNgx010ndFh2UdsniEWoZ+Rt/UclnV3
F+IT9cjJK+5T7UR7yoyyxzJhS+/V24+ufqa7wpisdIUmeyb6ZgXkCoJqJQinFDnL
MedAgFktWaDxhcYigViDgsWUpxZJD5S0w3/riWitne8EJ3GxGpD+kvpVDhPCns6/
PqL4qbPesNHHCaXWknbpWCXTe0UhQXFQBCysR/18ACE27y1b8rE/nmfVVkMQGTLp
Idn6jPtQ7qzzNb/KlwPfCsvc0+ktFOKtpHeYKoUsUjYpkfB6cbN+snQT42VBIh84
qRyF9LGeT6PY6VeyHkO9LoBHCaWAEDQp0hHuRtgm+9oM1SoiFqKMnTKU/VMlsoVM
lnfcCiooHeIi7hh0/fPXYH2qoNaxNt2Ce+0sBwaSgArm9NsZP2K0FFok1DqZ8hW5
vqqm3d4vqMCmNE3A6qEWGE3/jRDGchZGxvd2cmvwfjQVPfOP9/v0ZNKlsXQWLeFW
/bSn/RQ+1AMxxbgDm8paeN/aUfedH/XvtF9ShMXDqZAsSr4dBhfIWgBzp7OYOn+i
URjynA4OhFh1Qs9lpQ1dqVUUEPCP+MSraZm7s+nPfNzNb1YP7En9gbqloZOYbY/a
PDTmX6DLr7MJfCXDH4e+tK4yT9eXvOG9sk65Ud1y6FTzKuGsRgWdnyfzLz+dWL7b
jo662lu/Fwm+7TLtKK8J+1LYdOQTNqKEgCVQV3f7NA34iTbkhIIFG5bn6LEHeDn0
QgCpwse5PQFVXbD+vKvFWFZjmIz/W8oDNbV0hw7L5mGIk8HiSA/cN68K3hhWN5SI
X+hAGOJZD4Y0pQ00VDNLS0F9llps9yaE5hoqCuidh8N6UiK9FlaBL+dfm+UA3oDt
EOSRpK0/MAJoSAHmp1BUeQXOzmu72ZmNcw1NIcqg4MLyV/A3kioVUG+UWXCsF++k
tHBy/uGLALlf0+TTIRmBX0X7wFFZd2j8tMPjLn+TrZMeCHacCb5d/MdzG+9myjds
5BFPv0PGUYLoUNXnvE6k+NQLaD1/9qj4vbJxHo7tF9RBJLCyWmfJoB2nD+j1Bu1T
QF3UAVj8lIy1lWDYAyzv7yXIX+9MWlCsuHsclhKClGtTrpQP9xoLEOIV0wMMEJMz
L2diUn+sPeW2J5Aty+VtlE3CdU6/xhYcR1ed839iMMQCBUdWNEjx9umuWPjqhQ9k
dw7/+OmdMJt/elTGmcmXvqSlGV0NAaAmhPZhCJRD0XxE6NMYH6qDcaXnrjxiHuy3
vf+byLew5mUZZ1DYZSrDVhbvby8/U1FJwwZ+wWN7KOyU1+jiw2fbsX4ZBZzkxgE6
+NVBfT8tUAIABecnYMvS/Cex4ZdGx926uLV+zrUwWZKKah9sGs7SFrwPzXPTeXMD
i93EhAGi04xD5m0Ljmu+5SN7U5Qoa2qKn+i19+daoZ6GYjiv2IG4X7Jn+aAdfUOF
saIhlkVusZddy2miQhnkqcLQTxfpq/rYD2lACHPaR90bN/KFn1ytNzJxNchgpRld
0a7w+0Lw+JgYXvibzChizwiQxeCiflU+fGxxb2yVu34TcLW45mUDsPxPRItroqkW
FwSJrV2m37H7ajNhAPblkl+0UyfJKSZzQWN4+Vl+cHajghwc1szPxKnDvF4j4mcs
nTP/h/GhOdZM/ooGRUDA1QEYSfz+pZekFtJBlyid8LgmwRm8epCJRuBs4aNeBkdI
p3c2MKYPo6jI9BXmlv7A4kJ+Zq06Gbz62DM5GFFLPtgQGaJJKdf/FnCJ7iExmFwp
QCiNbknfyB6j8eVzLcClTVysAHdIL6YsjXrkkakFJMumlxmh1ZAImmvtoOF6aYwu
tsngc+wb5iIR4oP+FiggXqyaVAULaHMj2iZhQZyvzx462NOuDj14Mwb46D4P5f+R
E+7xcRphdCq4BZHz5mLte6MwBwcASG8J9hClqzsxGt34gBosYJrnHZY+1Uz0oMI2
TR+Cybl9X6Yf9jPyTh56QflhBiYJSQGyR5fp3Zfg5JPHY/gAn9I3uB7WEUo67snr
z79E70mrFdKUhKkeMP73+foVIcB3Oha4k5gAwFszgizrH5IF2iiCbVN59VlS+Kss
Op7x8t5qvfitUe9ZF6/TWJS8YyTNQ5B5kcXjBVeZJii74Fio8h4VBZWuPdGi/Ryc
9/8qyh6HGFJPs7HRXH07NtVn5IUZ6vePriDjLnsyEFJVeNFw+gnv4rO2UkYjOWiv
0wEC6/iUX7f1nM+PplZ04WstQhePwKTP66BCDiQkkfi92fo9J6yhv19hqxBrkLzz
nv7xiIZHsawawwcWwNm7nWhsm0Pztk6Pqi0frO0Y7vnjCjr573PICJCEq7grpKc/
bfSJgWuKwPZijTkkyY+/I0feg+yoAKkIoafjAqh0AeN8R4Tslec2id6VBxehuka9
SAr4gCB1kPxm1jM4jRBP+FYbV88R2GVKTY0qCXK8scsj9jVagjo57OPzKUrRaeWK
7BGFxiOWUOCir3K/ljhiCDpyrzGhQi4ZMWmHTsCZuUys++jmu6D8mRGZy4aGG7wn
jsA3Vl4VUq2Kh3AxPxlEfIiB0BjhO+8x0Dc8pg8Y8SqGByt8uVZqb7j1nEeAQI3u
9BZgI1CzvZ44qFVYb/vxHAfHFsAJSDfhRwn9dI2asJ2l9CYiN94HVKb2UsuE8Fxj
J8C48sNhAeCy5Bc7a4L4SHy+xImb+tqNrhfAaCuUXZKuTmI7fkoQbghPfkuvG6l7
S+FxOvfdhy7iOtNR9MvTvVrCX3qN3kLLU52Chsp21X3RH6GiBw8K2g0PpU/WD4Hh
r78dRzvyrN4HdCxiwHHrwxLbDDAdyxFTtnf19Up5R1wCQ+IOB+Q+C1zMNLN/em/1
0ztclEsF0Q/o4z99QgojuydEfwOwck4iekpALYCOT0gkUW6ZdhHW7+MkX5vJJks1
cVlNyEgv92diiTd/rXnLNYNA5XZw9Qk3AkUQzpKG57TYcOiUZz6DV7Fa3gTzG2ZV
5zQ62yt5n5ioDjWj93NaHt/WiRk1NWQ5TYG/9IEONgQ0QVO1HhyzkxViwaXR+o+R
2x38Njt+Ptj7GW9erxiePEmiPxE4no84MD17np2ynwHPJdvIea6oxDXVthLxls5P
YiOgOwsgUX3C+wlxrF6Dq8gOVJa0s9iaSZGyZa/UuilYg9MZTwPMRhDeJZOZVS9H
Bcur/fCuhQaWS3ldGyZcIh4JFJCPBAJzCny6Do2gpqQ9GQDGiLnSP+y9Orq0ju/b
S5JML40acdCAaLJOukwTXY9iM4tHk4gC280fxZF4JtXnj67M7CdpLYf1iZGxfldD
1Gi9tWdOjfLQ4OGN0bf3UNQxmRnp7aUDeyr7ZxahiOUjEfokX6ZJuWfYbQePo7gy
J7/IovZ4y1fb6efFgPvPnLbXXIUn7iS7c4V47ZLcsdX8AK+StWHBZ/xn/T+shfup
1hPuI/pCeUxaBPD443IsxRP93G9t/b/i8EldZJEiCHMW9HyppnXNPy0jK/CYeppk
TSZ0BkrBr8PHqF7oCRtGOyyLWgHA7zb4G3hmYuCtRP+REKGbimroymHvMRF55ymF
16Ix4ITMi1V2hdA6sw4wYwceEJCpj5zrguxMv8CWeP1zaF2S4cOGkf3pRJB4HB5j
daSyhUNWEryzPLnL5ADYgmOST8jJ3E+OaHoWenKt6qiORcS6CMq5LAiAi6keUOcI
CAu24PUC7PLLuVUKOD8TDtUdOQ2OiPJLaIaomC0zZhYyZLrrH1OwhcDBg0Dg6ZLV
VGZMxjYD/yrgYvA9Xf+Rqe1Z+Fb6sjNpfpqOnbuBN0d1YOTEO3rIF+nfL5HdAU9J
paqEp8KlMuYh/N1BE63S2Q9osxHrD+egq0d2xGqrx17NsvQMPwM0gQ3MoIKyJErW
kv5UQfjNVo3O7mIP6RMyN/F/0FNs+iYC4Q8cWKE7a9RGcukjeLmAiRhh5z6qDcob
VT0GCkr9GxRXO100ESGwT1Z/6JnokJhOdNWCtyhT8QLjzZp6mJ/sSQKWi7kRVKh8
zcvt50kO70DaFy32149D8/e/imBODgQoIBJvLQvAdMdZ9bk8wCYe9si881OB98dY
JNCwCpF71LV6OjDAXtAKXA6cf23cjGLlA4p4HDfhgmodLuQg4NzyQrc3SS5diATQ
77NhhF42Q+H9KiL5NLgFZu0eud43P1Dzdc+SFiXyuQBYtvNQs7yLEjeWtBOasNGD
E8rBfzR9+qvvFCbhkS9CdznMrwmAlVMPRuY8FctaMsmMt2lKxJRaq8JwG9zsVQbl
WMWS4TCr63WhrFQDyfIWlUwARjs/2pwgWAybPU+UuqdU9aQTBzhL8Apj0HtxINCY
bYWfXyfhTxIXYAaTDPN6tUJKyJrcG75IVvSdgqpAXHS38YXm2RQBYoSjKWp4uJ09
4dpMtIB0ahXihCchkEYZgoK9DeHjclOmMMFZk9SFKjuESpkzbaF+uAWeXpTCdlKw
vZgNVTtgH2Gru1Bt9H+wtv5cWq1qrfIeJb8h+u/xvCjyBiNWWbowpEHlRpbt79y9
m4lOXlc20m1vV/Ad3GHR0l6xosTyFs4mTpCwwI8/8Bx6NYY2pawNJmMOuldVKSEC
rTjvOvAjKLPqYhajDPbeRTuya0Dq/JI+B9ArJX1YNMBzhV6itQ90tWVizzaZHfNi
hOY2GO5nZpXs46tcT8OZ6l7G3Ba/dDIwojg5Kp0jTnqOY83dFTLWfDLgUH03owTr
iJhKt+GegfyknugNoj0QgSiwgX1kzYaicAP8Fx1lTu08F9iz7nrZNqtUrKwrigsV
++Jn8/a3JT7+U0EupxfuxAmtj40UkLVc2pOYDmAJCIB0kRjotxZ+c7rsWpqm5ctB
QILAAlZE9LWpD6h/3d7OHfc+Erb8oRTua0s2/SiyS0fuquaaGtWxh43voEGPeZ9Z
/3eXwrA4iAdYPeuLEFZyzMT9ILhmceQdLjqwOaKB9m0AnY1Vt0/XuNpjis0IzAF+
aWIPdeKe/Qis60etxvMN/OrnuYo6Phy4HPMK/j6+TGJoyvrNO85090++08Mny4lu
LTOvwZ+IHwreZC/AWJxMEA03k1Fa+qWJXlYFVXbGnQjbt6D8MywR6sLPDgGFY/zj
kXkl3W+WVaB2gbczCkYDPNgC/IH+BwWbUaESeKo9dx/iMumSBZzaDRVVJ8EQeTyC
kZu4kuzfEufrZGUtgQn1+hsTcKE1+/Up0ain4d/QTBfFWBWuL+j4KDinqLAg1rG0
NF+yB9dxi8E1hKSc6pphQEGhGnGjNMNXSmeWu7uDXp38ozmBlQUbWFWYGRzahuiI
IonGQSgfIpCnc3dISdUOOQhyiC5QycZCCCTiagm7TeGsKrmI9a2bQhotvPymLQtk
Ik0Wci5lkUCOMxF7j3MPQaOBZIjNkjK6NYNoLFUFntqhN764I83KX/T2IdyU0tle
nmmp3tFJOLTtruHm92NQcpyiGagffUQowL9ot9CrX24PLkQ3K6DMP//xhVJG46wq
h5S5Jrw51p+74VDCpZb41wI+ElfvdBsqSNkD80DdRqI=
`protect END_PROTECTED
