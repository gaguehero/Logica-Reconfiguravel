`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IvZLbYJ6NyD0lA7RqmbSRphBoIUIiC5VXRrDc9FLh3SR5VM7BEIReJJNKZSAYwx8
Q3X7FahzrCyR9liijqZeQR5g3SipvG4f/Vi8iPzcwUkvdIXuvwl4U9U7VZeldHLI
qIJNCG6yPjiso51gVn5i097vXb4G6/qJxy2wuf15Ml8yQtvMP8NPFMlQI2M2snms
vDiuI+2g/ZRFw2bf7jEuPqe/wbaT7hMiaNpc/NbKNsEtu8uWTVJgavJNF5wj6F4E
jQV2Ivsi2BycaV7rthd4prAmo9VTxAKL3/wLr6HhjeAmorifrHg87VLDf124OZYp
uXVrhduryI2E/R+uigkhEf0D1PFO+nP8TVny1+zR7skFwMmJhFHSqtFUJ0nXVZrN
UB5aFqZf6EOZtWxpoBk4zhNYNPGiFfR7vrBm/mfCTsoqWVvHjcBS/7t++jl6Iy+x
sdANphM/6g3wJHLu6DbEBULSPF0n9WJRIZiHOiQM37uucfst9vH+gXVxlPfu3bPz
tWJKJFWBnnnq9uMKdkR9ShiwVJwdziT5gcHtK4t9HbuHGDsHGcquD75tHp2oX/Lh
fJ/KorDChYoLB1A94igDsfzignO5WkiHg+f4jxOUwgAoA7o/dg1XCEaPAev+zwjV
ynwwxNtksTpJTz/yVuIf9UA5jwgPkpd2H/XLn3lUGGWva3wAKF7dA0S1018NYaEe
8sM+md+uTwSORo+KM6RtHcFm9fWfHU7HbUmB/Dm3TVWSUp0rMHR1Ehi+mm+wH/pg
y8vPzbdSpRwfzQfbqebp60XAZi6Wz7liGhq7jNeHGh2ZS19eQBcpW71TW6ynAga7
2wcvRaKpt/McFBoPCJGwPOIPJNULejvxT6uhzZWlJuMB7LehBvrIro130/pyD+4P
BQIbTnsooebq2uuU7rMhLMkJ2gm2HsWfynWGiELHbViE25JIIlYI0h8egpklpVNW
sCIrL5JVblaXj5xSwqp7g+qnrHKXolEx9fxtQAQQtivprbPCEm3Dg6VVM1fYRyd4
HGPODowFc2Xd3iC5TCmnVmuO9ENhssuN1aVY5vM81kmS6Y6vFf7Q+HRuUw/U3sey
pOjOg299CvmNGRmkEFBrg4SQRx8D/JHHqPa6H+Olrz7X/56SfNvP60ZaYs0uAiGf
Q1djI5Xf6yyyHwwdTMINRUi0Xrt9N/9o5TokjzYHPtvLmWDHKZy30KO5XpL1DYJ8
iqPSMb+Yyplm4Gew/cMjYhqUMQkbaL05Z/gXM41/SXfCVjCt2nuNcSK4MWRpCAq8
ZGGsgw8lBg6MZUE8TaTF/4CCyfedk2hL//BtoJUhlkiogAiX4CtbsYqLLNFCvVTc
x0SftPFwhFPPi7GGIvfam/d61cjFKL1oy/8V845Qv1FVPOELF2hsn0PUeKaeJRZQ
jF0Ij+pJTGagOIfj8K7kDMc0lLsSOKoUihjalYD76+UHbElKViBIlWJOTto4V+sq
lmYE55lLhVMwrUIbd8i1qH7CzbvH58UsVGuzwVcio2oHMtGdXGyvGvc818abRBzT
/ktmWUNdmbT65h5GdGqBhJ5TAtQ3q4Ii6ikk7IoGGvUp1qnFACc5KXg4y49o1aqW
OKwWIt8Vsv7UUpKaa+/DqMXSpbcN/Yimq+vZJVPJpt1PfH7mLxX+7YPQouEIQ7rN
txSeASbxTpHYR7Klzx7OazFBVAqT/qpWtiv6YzT0ia+PwA62xpR6/g+x0/1TxNwj
LHrEnqc6Z8fDpHS84Tjc13zeWiUzjGvbI62wku0IrtNZ/zJxFMqZVk2/ehORhlad
uUcsteLycBYjnYLMnkLMgoR2UyO/7eOE9wQFUke0jjZlWY9U3Pis05XM+DUw189Z
7q1uX942OtKryitkIKa9zPbSdpEu7sp/CwbKbq45i0f7Llu3ZBFqupolwSVb2R1C
rquWC8T85B4I0ydUorEYntKp6XRFJt6uWnp/xIsq7T3gv4TEnaWxdYsZCWVqOLxR
Kss/F4XMHgWRINW2BAG1VuMp3xeLOqHItDUw2ggyXX2Rjw7g+heFMDWArH6mBKy2
yoarad4ECogK+FFUAkaPGL1BcQUC0mZUmzC3orRVXTzUUFBBocU186Q3B34A3MDd
lrhVgrdFf2sT+w0gzNG+ttZnyjTSG9iG877XWUVHhAuPNFOyraV5fDGk0IWM1M/h
nUXUVxS/VQN4ezWHfiCg3zu8Sds1oJoYPxvMY0amkNJ7uoeBFX+E9bAFAex+aeLn
xQO0W+o3+4ZFPP4na8B6HQ==
`protect END_PROTECTED
