`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bpQgB8r96hNyunM7fZTsErS5Cvi4CEhVG6wye14pSTEXlXYshsMmDyLGLJHckC6D
Xrzc748viVr+QucwxKXwFMfyCMYZUfik0oraGI5TrPp+h3mqVuJ/8pqHHu+iLc4H
cMtdF22YnM8VoROBZFixvWmqnqxDMlwyd+0oUz5figUiNF37w5r0tMNUanOeQEPU
kmIpuU/y8+qWUdqoAotbDEMhmX+mPoofPYUJOigLO6KiWG0g1csnYJiGIU+g+ACc
LbMELq73AI4mnJX/8ZOfxWSrU+mZQ30AioyCY3nau6YrjVWss8qOKo1Edhgv9w6D
6xkGQSbR2JKsjtHY3VKPavl+/GMBsArTO2YqoTDzI6xUqOGn1sanZmEVzN3HN9PK
dCOlHp1sJs28PI9SMIbrq/TKu2lHMXnkV5SeFXTcm5qJFkZ+GQEUzc+uBIrSLMiv
JjA6xMM8DR5k2QvRXbuIJX0r/P9GuwOm6irPZDRVIoDIrA/H1bbDfq+OLFGzxOhx
zli+/Lj0PgLnD34PNwx18jFeNzsVwwZjrHJn6kllr3AOvsxg7HYA6lBdWQ6SbdGo
ci+nfMlW7Gl0NOMYn2ewNvUJS1qZtTbNmxUbvoz9AHnFIul6mwQs8U7z/qDF1JLN
zTyopYsux1j0ghhgvFBRL0Di/0DQKoB0z2Hk7rEA7oMaiJox3W9X5uKIIbC9X6Xh
z2xYbWdRIa+mxLijKjeGeySOHGVK+EtZ45xHvbJ1hPMd3FGIieGqIdHisDlfmcej
O+bopAGJLx6vcwnoLKPIOrEZtxY5Vnhv24qmHP/n1R9n1yWuBXYJ7aYxOQlUASis
fxGNLBAgpqGIaNXVJrGtK3vS1eobcaILHe1Pwe0w8hdBK19NHr1ArFUySHM3v9pr
W0Lnqn/nXuP2VmqpKesmjfHDhD1XcRhjZG8kmOSj2BvCLg7Fzm4lS5aXV9EDV/GZ
xo6AWCA+A4tUcSwfA95y8qpGqhsABPI39SyFoh5uxnp2gkQQR00sjW8xTuKW+MPR
sTEkQIgtPMcDThRoHyOZKv1vEoUir2FmcwtYsy1sqzpH1qBbaxWoAwm5Qjz4GF4I
FWXA3jvxGXTmv9Nl3joLM+GZpb/uBMBpZ5w6eJbBXZECxMtvKLgQ1+gkKrpGeg5+
6/E9RgPvKRHm34W/9SQvTmiFCFuOgp6wdyVFLcCbjEDc3QfGZKlzU+90CJN+PgNd
dNTbZxadHlLElk4v5BGKtTgeGUu5+p7V+v5LrRAnqU5TLprbNncjMizu3NzjUA8/
GuxTv60D/e2/K/weu3IdolM3MyGxK3YfMineSMDrIntlPaR0A/0v7XayL1NMRHPM
Ck0CfqJ1mJKq6U83qT8oMYwLyM81J7eV5umSEvBcBVbSFxkrfM9Q5rEedGwwLxIW
JZJ4URoOAsDY11CbtD+N7sGcODEJTiWl5UkQNKmWVEVihT96g/ymYdfDlr/dZlgk
Kvx3UCww1Co5kMCjkRB1Bwu8ahLPg7fSb5bESF4Q3AS7Q1x6SFbtP1kt994p8gFj
O+IvcmRmxnO7+PNlxrEQQU1Cye/UW3Fk6DFjLDQBdkkYOV5scIpKRP5yR6P/R4tW
It1WzQ11ZdCgq3dj6JD4JS8+sL64FQgedc0cjpUAeWIx77nWYHD9A6QiCywxNwOa
rEUphAJt/jBrPzw/3Wza57t1zvKSN+LI8YbZDZ/Cbc7JTrCRXvrto2jrDpRj1iAW
8LcjNxBJSwcRbz5iTvrICM1mdY+ZJhixfUiw1//SUJYtd0GF+PHRbBN+EynRT2qP
qeK/wV0L/omoDtQy34DGXtc6kg7oiZ2mkroF4n7/Eqv+jK8VSeG1+NyWyqW2gt7m
Gb0V5NK5mzCUn8ZG7UO/Kh1CdWeSF8T/9mFT0mMDhj9bfWbEHDZ5qsLqL+4kot07
iRXY4lB6iu9knitHbaA9t2edcsyOVsipe4/jEd19/7Vll21N27yUySo/+t/wFm0K
fbJhoA1ubivvqBsBDe1boTW5y53cwSnhp3xR+YxWI1C4XZrN06faGGNo/FxRzdvT
6Ls23xdHoRVFe+DQSBCFDIT1cLF+QIe7kjLEQmZV0DRuIAKGEAOrNC5UA4Pmff4G
dk7jmz+Po3kX2PASVgcKcgWipXnslkg2eu+IOx+hXvSjetL9Z/DebjUF6AWNbh4F
kIHF4xwI3SsVzE/7aIPVq+BdvrEMP/EVUDMMUNPCXxd6vS8I1OMLV+slIm24QXiE
dfEBG73lHiDkd3NX4j32W7/rPmXXRoFWVRgtKnZxhOhVN1GxWpBML5eqyi5r+Xog
79IwHfw+P+cup4B+L0dk4Hl4qR7zfviOZFCYE3w5O51P9sWzZXI0p/X2dR5tA16G
akuh/C9xLrNIpGkGxR3rfRIsfZ6CDJYAEZO2ntg7EX4rS1v9RN9HVYvQTq+2sVcS
usrXVqgx7Xwj5Y82H50KIG/BdTG4jan3DD4K3u9gtOgTwUzh4M2jizTnz4i4/xEE
WQA7prB4EczJ+XCZDwM2FxtdHk6lZq/7A8KlpqzZ84QjiRoY3O+KYihze8JbXbqo
2GJs/khxTBBOqiZu6HgPrIqtgvVSDM6trMNkICu4ZHYf/50frOpGYiMiQGC8QeyP
6voDqLmFcsHxwrieyjhDCiQbWO+rykTj1zvIStWiIXN/KViPCARu06S8QK39aCbW
T5cttr5navIb1k6tzuV8wx/1adAZh2lmsBSx/IlNd791XP9CPRr9uaJc2ejLDMrD
BqNJoUg/YYq95oTHgigl+/YicSqiduKPRPyIUx1qbxQG9W2n/AsJMjdQgeHhVrcq
vYWc/1cGHakG9r7V7p60mDiyvQIrsVeOHkPL1jm6/+NbFwYexGzJqrrmAlnqJ5CT
Vu5pYY2/faIAVnx0HOYHf7HbPErA2WytvJBwXX47KV3lErZTroWMuX5lZhtvd7xa
PG8JyMcM5GUlWWKGaV/88efCgLLJ+lJB7p315/Ew8gjCfwCghsTpUR45eiNBHVG4
4zrSp8/vyiSX4eSlvawW72tc8GGYBsC4R+4Srdq/ofKBNAr6FrwDp2+uzVu43DUO
bjUjC1drDOmnmmvZJ9/4o8FQREtBcVEMBdGmc9nQp/lWKwtrD+mQrYB02PNtKRWg
js3rUHa0rw3zXR94qKAiCqkEWslLnHIFExjgXuYJHFURi33k2DGCDpTAVr7AxnBb
pvxa6KfeYGjknz24Rsfvb2N/cYmPcW5mHu6PXkVKA78de9ETQMf+ipbzrvkKYi4p
yGT+db2KL7G9C/VZygqGlGDKj6VhRXrgHThcB9e2Z5ATIOu+nIn88gmp8exDvNXa
aPrrhAe8uHhRdOc+QUPJXAuigzOgvPQgwlKV4Nvi7Jq31SXCOhRm/CIW+GsFApN2
63IM7V4f5QIBSgOS1Vnuj6Z5spS3+0abCWYoC+/ngpa32Eebwr5YDWlJxmFfslv3
ch8weelF3oBjEoApEHq4gA54zuTJzsxKFTVFDt6/dq1WZBQIZx6s+j3JQSIW6WOU
68mO3baU8M+wPJ8NpBEezrKb8bsdl1C/enUJ2LF/mi8/ckrQccQb2beDIkrvtcjL
R/dKn3GjFCFn8AX55GrJc2WVLkEG6CHJMusGJ94IlwCJMGW6/C9/dvW2FGYDeDIF
k+ckj1IoiWoVoVcFsAREIK15IUVyoKTyzpjO1C89ZCEYBBOU8s0d4aYcNUcv0ZUm
2P/sEkfUP/5t75yLZDhNUtBzsjXCSjEK4sbUJ/M3UeZdAP+IntVsXCFKKQZ8YswK
EZ6oTNafjpWI1a1i8+pT/JzRQoMSUUyMu0wctyoJSc4IZpDoDcvIUlBe+Q4YJPkc
Jo1Sg3SWymFTacbZKRW+SGvlWNnSWCRmt0Vf81xOyU+KOMePjUR4/FmiahTZ2iMd
4iVFOcV1tvMwywEr/UOLtTAloQ1FhDmPAJ0F6emWutl+q2S2CbTBpGfTraXoWnk8
RYRwh7o33Cp0W57gL7IHxYK/1rcvd+gk2s36PR77vPy6DANWTXRXs33/Ui/ZFBze
nd27IfFSTFDF3RON+WbUwsavUI1aWDW5eoLiU3VeuvJQr/gZwBJOwBZQ7HoZm0na
qD7jt6Xwa95z0qfO4iwR7DVdAk8HviZ6DM4KeW7/3j66qjafm3NcGPW6AYrbUKlz
1ogFkROdJbj3YzOyRnrqLit+UwfsK6xYawqMaQ7VWJEiLwUFGv4LnsjnO6O9MbXr
NRdHQGKcWk4XHcyTHTsLwm/a73qZg4+GLa6NrL2jNMUuBMR0EB65kmFf0J1Cc0XB
tXFHen9DQj5UPt/p/Kyfz1WtMlyCphnk0UmcpWzz/tBxjuPFw1GvvGJ7AIuUHF7V
I2gycn6RB2epgWJ6gxLuV7EO9vOCJsAMNAbt4TcAK+tPlcaxmwD8AC5fN3VfKioT
AzncJEAGcWiJQ3LHjqoP9xJwUJLLgU7Ucf04tyBPbECBQryRV9XJg54i7lSMCeNK
BTgmYOolCpieQ6WVCmr1mRRKjJccPfBYtx/B8Qz+NUlTNoBVZxbaAAlrfmviRxt5
yHVsoOv1YaKRP3s4vd39p01M0nuUk8EohCY2fm0+uzQ0FIduZKRczSTdTDNacT/M
I6rz4uh7XF5EpOjfbkYY3RezVIcSLRq/YT4cfNwmcDkeeFCRTxVUbgJnPPzc0qUG
Rf3Y8nemsoRoDL9Wzv8ewyEj46ygfYOTyCg8nzJ268OY6epxK4gP4MYIG31EsdYm
qju4sg38sqOgtdw7lgMRt6fG5ClUf14ulEojG4yL8K7u1fhC8YkG0OQMmayazrEY
ljnerdiuWn0tFbcRfLyt4amRFpeRjU9i9CTFdOnshNswAhcRYzv4xPduqiUITr/w
kHLmkhDQvv57EMB5R7Iy59XETV6CmbkciD2iZ+ZnWC0W5lJfFRDS2EmmQZrbwtp2
4esz/PeG0CkquZq0yyRXx9JuMdcarNsFgp1XaNKpj47ZWRus9B4sCxl76GCQpmYy
rJAcS+swblZlmpyJSkQ7RLlF7jYnAVAU3PEYrBJoW1CnkwhEVC6L+t7KHugjzJgR
3hhAoegWKTGtf3TWEWtjKllL49i6KARckn9gRMCqRtFzwvXO908HuRdyF3Uwy5Qm
YOK6+K2Dgl9O0hpT0Eo1lnL8Mr+8NIPK13dlFAricvtTbjperfIg7Kts3suM29wh
IxzDi/V63yg+3XtrX7SGDe+yYxs8phhOUkvkBri+zMqZLziEaKkQe4OYBiuhiiu9
TI0xDE6dimfNoLO/DDLVmIVKAja1uQCQ4lL5sJs53iOlrU74bhNt7zmgaAVBHAwA
LzTVJBT0fVAmSaEcXr7uh6JMDI6riStxymTcn0tcaJJtrCtcXgqIU9Gz7Ha0ZQAq
SG1TOdIYk8B7u7oUmd30/xJBG2bH9cqCB/qB0LIPARVS/UUdrcjsVkY7+aL+6+Sq
Zb7XlPvrKVxglfLN63RIMSccsoQCAjtRlOTcjDx/W1cUqilPxkk3gWEeODBNwpwJ
cfdX4EKjoU8hs7Mwf7nHhg==
`protect END_PROTECTED
