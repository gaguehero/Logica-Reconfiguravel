`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z41zC1JeaZ4JIHskjWbMbd8UbV0qcG/T09+jTaIpEWT2MzXFgA2mpffudPG8et9f
rCy6jcK1a91l/uQnSTNs47oCLdt5GH+jlz2SGSw+vF6hZ3y93LOdd6r2RtP05HYG
bNwjKBeZzPF+E6EKOnyNRo/1ZoAwgR3qyE7KKXlDKX9YIaXOId5+vDdrjCQrjFW1
kT53kr4oqsGZ9HDxLgiWum90KGyIY+d9flM+fVqSXgMQVfo5UuXBcJY5gGJjpnoB
wQ+yyH1Ur31E5tPBvPts3qX4a7MX01dOlMpsohWZFWQlYFPwef1LMESIwJKix+r2
TJ8vPeTZgzzdkeji8Dd0IWn7XM7ALlzTiZ3UkHMFsKUoWnAFoOuCudbsJa0GABL8
ID2NeCj6yhDQWe2Y6mvTOSzsUjwDUKyXkKVlxny2M6fnD3afVxkLDlh5h/V5qED/
siIo/PuONDiw2294vcrOmAfgHt5BeN3rxlLTw8U3aHTl1ngU8RrkWt5Eo89n7bF0
dNppfE2LqwSUJyNYCfbHZKnjlheUC9JkuApuUoZkIoC/eFD08OApFv7zoafYVtaZ
Nvt90t/5G3r1yJVggQJCl6wL/ZDQoeyjzJhGLclVodMvLhut//WBZjSHTuA5GT3g
mjNKrhY1V5LesYOZqkhc5BLsALWvpn7GnhNuHfvb2z0EcfQer0mvsVgwnRnhPKDt
vxFTpIPBZve1fv9gwtoXZq/863JX1moCqWzG682lTEPBrl9Dk2pfEgvtMfZdui5X
V+lr6gbpXn/sGTfMYHt7lvtx95vnSpWd2mr71Sf8edq1Nd7zNkMiDUq4fjwwxRwe
vaQ8xoZd+6d/GqPEBXCCBP57BUD6c0MSepstnQPTsoRVxQD8oCa9Q3fjIHxpbwbf
kykYTvuVoYNDM44UrNGmPfeo1INBiJJKwNm8SSmgpM5uMby7FwLPKahDsPfRjoaq
CUvsAr5ADGwJel3EdMpI6OJ5zYdgxCS3QYdiW/lKtzM7wSfQ0ftI4HBvOTnYjDMV
E/wvhvYwvOtrolR+x31cgnpg5oy4ylH0WALdHF9BEPv+Bfzynzq3AEGlymANx01x
YuLU3xdYtk1u+nhLPiorMAaqOpVT25lHEyeUzQCPW2K1wB5ii6yM6GLjknoR3TZi
PcjmVVM+/QlZ/eDuPJHSRu5Rcnds66zT5cgfDZkaHZcySwyHyk5RevjvKGITSiQw
KmAQjfS3DfCh1Yz7mKGxJY2ZsjiPtpcq66brvsVEKbNH6YYKI5z8VKjfAwNvjY/O
mWBn0XDDuUYAnSnn0HHH1p68+Sp9GvdzHo9TwLH75PvQew9NeEqf5K0wAxoiMWCr
drr1WCgUQ+tO1XW3kRsVFOnY76Zd4gF3OXbXeMwNo40sA1kQYu4twLYa9TxWZjBD
xN7ZQhwVqKtBot2rEpogzG+G07NzdsDu5ZG4o6OUCxdpSxEG/eMH+thdL7ZX3k9f
sVBt9oz8fSF4cJI1al7XGVEDx5D9OsWGa5wQLBBYiqrFa1slG0rqbiiS8LGfqj4e
GLUk4mKKern9C0e0N7wQa6ZC+ZBZ8VLbHvbGzvwsNbd5wnCoggLAZ8rWN9bmNMaE
RaUjFlSw+CThwnxC3CEU0oDiWbzu3vUoSVul/EH9AFE3jeZJTAB6hRRzs8BSJB4/
jN2DKXexgIsnRjNCliyJB81lnvV8ryUhHYLY0J2KgJPbbR8QwiBSxVE2vkHZcckc
Wp3954yoBe2MO6FvkEzNfRgLw4cX2jYSPNsou1OoBwBhhRBZwBE4DDP+eE07KckM
PZe7ZyJpEzK7UhoQnIhoyS5lIU+CULBNcP8zqhUhi5KgRq4hZVyEjsiugXc1Nl6g
Hox+C+LpIMVuW9j8s+9WwGv6Zt2dsCsmu48+dixw7wnluojEW19W88hmcfeJvPud
Y2jm8Xlh5vB5UiF54Q2oUgmwzlMWryZQXJKkt5rD3XF2G0tHHN3OuMIA8OStc1gY
7N/VCQEx+ZkrGXTqQwrzunpApG9GVGBBxE9jhyo4oPT56jUbUwtLgZiwWDI0lRK/
RPsn7eOk2lx6BhDHY5TgVSStgrLY6zbU5/zrCU6cllsHWIGb6Vlrc359vITkgZ7e
FrwyNY4N9D4o5KQZpLLUOOHf7Bxzyq+OX1iE65hnKFkr/xgpKaQp4wdrtFOTnoJj
5lazwlA91RzhpddssfQFqgfw7DzHFXPQGKrH387/GTrXSX0Yt6haRygN5wW+yong
8eYwuMD/q36KahdheETjrQ==
`protect END_PROTECTED
