`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRa2zBOGJnNOiiGRHklhPxVT8M2fAzgxobK1Z9sqbO/Q29wcNyxWqIA5sZtpCjny
BGFWQr2rGU118UVtbGoEHLtUNdcNjhPE0RVE/JGSpLf/HciCJafCbo2r25uaERow
CBdOmvJCeVyPt0g2FPBfGVrlK1e7fjz/Hxyf0YZQP2cIwruFWPsi6TdooYgCB558
B5O+8QPFroJGC74L4d3+JGHlVl6XvmJ1/GxDv71woMtoVQJhRowFe3CV4Ww1EC35
yuEsPm6nbxrGQ44QbfUV6Pk2bmTYbF4TkN5+Gj8RajyLIyh5+PJykIXfs+Z/t9rk
k9p5wDAUHkwSAsdDk3Nc91EkfhCo9lAOck0f7iRWoCdxxqZAEIi51WUWd/BaFtjg
5J5V40X59bhQyj+W9KeQMkX8frnMzkQ2DYDDz7aexI1TQXnWOtUXr3HbvFerbYs2
Al9qcsvN4x1hQe0ib5zwfQ4c/gbRiui1wylKVNEecr94jVcTR/s6ceDJ+hfPhGz3
8nKijgGtnaSdby6tCZp8Njo2cuemkEoCXwDo8u2MKPFhsTU1xhay/Ud8pffnjItO
eZuwl6Q8thewdqwXVUMfNieEpE4xyBRf7E7VW5EPVuIuAyy9PDCX8PEVZPfdIXJ5
7i24ocUYImlc/kLPY7wC4w==
`protect END_PROTECTED
