`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4lkVZmLspsHz3jNsYkmaw8uDuWPP6Bcd2Wr9L7jn/JdJp2iDu65mcw3m3bwbgdUP
3PnheVO1+W9V9w5/kdWjNmMEq2iYOsC/IGKxon6yQWLrXZZD7bDlNRRfbAmtkGe0
WP+YzWy9i+U2Rc03KjvDXzJxbIIvQG8azB9KUqitgfo0PlbUDfA+db3ruDnzfD1T
dy1c8MJTWvq7G/0wm/0GRB6h92OodBcTHD0hpQUkbLJZu8CgR3fuUJmMaDkjk6Cw
bUuuwHBQtC9I3tGFym7v3JwIDes9udEn5ckqfrpTtV/xgcu1TgEttv3+YIU+qI2L
CoxTRoo30Y/EfT5c/MeetmX02r4ppuEx1OepVel+Mg0pt0B+O43ws2sfTA4vmmQm
c0spNoqWvIKRJ7LTQLJR+cs/iRIaOD8cLHKUfEfzdCINVr596cyAN63IRAkkDGrV
+NhInKfjU+e7UukXFo09DOekqGSTDIkumedMu3bYtFxEtfss61TW6Tif7y5GnnnF
cAkbKFvowrOspOwsPPTT7yYmVUyLC4xb0RAnX5bg77HVG3hPow4czuuSH2qZEEAm
NB1DRsNwHJ1oFFQq5lELs1ZhABUZuzSPE2h7EK/06HOhbVEXJV8O6uz4xruQCVOn
YMSrLM5zHrwPUHCTkaep9lclSbaoB+UaAfRYxM4DkfhVOwQySf+R1TNPWXrO3sdK
R1xeA8L8LMAbAusLVvJIBpymuiHXqZ24QWqMi0vzGjPPy0Xotlfwd5TGz7mvWnlZ
OAxYT4ObL5smvP9t7hRtkuS2KyNzT3aT5HFmnT+3R7yv6H+TpGn8+TRHL3ZvDM9g
K72KCNCXfnHipe7QNDBbm9tZJLnsOaHDX3rYZskqMNfCGnZKDVp5IuAC/YFamDMB
vvbMALTklllS2H/yskfw2pbCcJqt5WEIyyai7BvNjN23ffAdxeDsnG38r9WQQ4DT
tEjTvK33KHUqBBwg0FZrkN+D36MOiLT/Tr/xAx9QqQrH0mXdzJRvpCaVMV+Lufv/
gC/3Sj6F+2/Ta+DlqEbzFng+DjmZCkvbPZXmttMMgnytC+sYULIvdjFFcgJtsJo8
berok82CJ2JrjZWKfNhyhNmeyOppME/mbtG9Bo9yNI37QqvhcnyfI8TxEtYV8Kpq
puwb+mdIfm8TkdOmiTPdDrJjEJcN8yAjk8PWfdr4V0nZOnyjJT8p/FzQr7eZ7HWh
clrl7wz3Wr08GHHc3xJsO/AgTeLb2dJMp4hH7lJOGf2VKzex6zMb+2r6nWn9wysf
3I810l690razR2hxSoxkUP5Nhu4Xhg091KZBobzU9FYTvMCNis8Um7o+9oxj5W3H
GUluLJ/8n9QhtCNp+VNVNMe+maWun2b5TiEPltnc0HeCCDFJoL/7gnIdiskW3Gyr
sd4rd80IvXhUhKBp8UJC8C858C43jarzb4WVdUqRAmEuH5H1W9knIYbVoGSrTZL9
LEkARj/7AVzK7yYciQUzZ+kEbX3SACV/votw84GyqzUmB2yweAh0rEUfBRaKKCqI
Jbya3GWBMbz3fPoav7e/mr8H7vKyFswVFehOsGoQ+g92aoMlSaa6ivbl8Vd3JKEH
LTSZ4QEZOC4Zbfxs6rsx8KOag9yqXM7OwJAkTUhePoK7Z601DgDBPI0QB0rUequV
Z/PAe4ohmP7ZOKHMXyuhPH0n5GDF7UCSIP8/NTmxi945coHjhDdOQmyMwf3W5XqK
o86JZNYICzAaWQemJUStWzKMQvZyB6N2H050W23G1GiHIUmVYaTQ/bQm1Suw3T0Y
8LYIjzIrfPuRRhx/zn6T1aAKCCSsvlVutX4ISz1FjNvDNpkUdlMxxNT05uf9AuDd
8eJCrAtZBmYxlTaAVBRjGnP0O06eOeA5ZcPLM2uNuFRNs+wNe2Ec6cfhe4Vl+eq1
7JoljF7zLpfJai3GKVX6Hn8BH9OunqmCDbyz/JuMcSXlQrISq5s5fchD+IRqVt7z
KVFvWuZo0gBG8r607vSNCS/e0mSV+hJbElyMHwb9PyykNK1n0dh/lRg2QRL+sFdx
ShiMHvFZtDV//PavW08PR4f2TtfS+XCineBDDE4qOwKwd84l7L/aILPh7TrbpQqQ
1/uwX/2P9hEYvYqUJ2wt/LQPrVCO5ujt5zPzOueqQFMILfD0KdRG6D895g7w+mFX
WNb9CyIUXhYh5jIg0zaibiLZD0UTP8JJiWAVrhb0OpJnC71YEzlxLqcQNNWi7Z4q
Mce0SNDzxxiPgehf3XYaNA==
`protect END_PROTECTED
