`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ6xanu6dPfN/cStXHgpfFmCx0Iz4V8h+lozVY1IznJzlpseLQUAMOlt4T8UuWaO
N3XYnB32K0ajhOO62lmwXoOreaQ2MLcaxToIRc3OvUYPfLKuZQVnfxbZS0p+chHZ
hmxaOYbiLPXU96T+kFiA/6In6aWLC3o+fSqYAhIUIFvz/naUz4RYEFbSVEgMsSzZ
x5zkGf88ORHEv3OHgFgwTuWQZcuAQPA3qeYUxzxGcdzaMNM7fiKiU8qA+e0kAunP
1ArjmLDvxDMm7mLh8nzJggWfUYAVl7Ymqw1Fy2W42zgR4V/IDxI/mQrlNjmNuPBY
FX282JkL4uMGtzTj0tKcFOlz9ZEy1pvHPu6TBLH/VEJr4pLxKUTxWHAGbVmzLjW9
49WsNvLS3bGt5UKNfv0A9mWFUoFu+XTn7FKfQqg4Vxg93VnWSaoXOwjbWROOJ3PQ
DA8eVqZe8f8XDcMLHZjJ3BkVT0NVWo1WvFYiJ8RFT1Pxo1n+Be2HkI3j5/lSv6kG
C2N07oA5nMaLqGtCCL+C3cVyvp2+6CmOIfqgwzn01UA4cbcfrz4L5GjslVlC/jsd
o/Nw7EmnWUMo8L4xytA21CxXULQa8HrQK+wZz42CdhGkAjGjwsXRlXWBRTEZEMZF
+wU1bC41lr+6Zi9Sn3KsHJTL865DyIxMJClWhI94UTRB8my949IrNJtPH0E1FqV+
JeqiKtmquJ7+nglntT1ue6HNwf/8Rfl3ctKdsTaCGEhtNiUxE1V8LMLYZtp3hjz5
exZXb1c7ig8seXGqL+zDJ1YbeA45nDH5a6Ckf4Bau4LHiinmvB5dmLDWyd28zKb4
3deKgKuibDk7Nril9kHdS8Da/WnaFJnyI5nHfSQpTVfrxbzRcHMEEXcgdhdW0rnS
hdbbws3Yk5by4wRSxShCFoKBObIcW0nWsLHOBuoht+VMV9E0K892wjCLJATt5842
lKd5LRljECusv4/0qmAScSfTAcYGWgHE/nJTnihPqXjcxjLhbsmuw1XiWs8Ex8xa
0ootc6pzGnq6gY7qPmRusWEsDr3MS9fzAixMtgNeYVDeO01pgBD2UVarOscyVhel
N9Vhl46FFVIcFonslAJmaSTnTSTlwN8nLH1yspm20DCfZj8UM6w0SW0Kj0xE14a0
KZCYMqRB66JoqYTPq5Ly5+tKMIGgYKpph7mVXRanzSk+BBzOTNXEuXwxye5/vVlD
+b95FRcPpcNZEyC/CPCMITl82Hf7uD5nJyUpPSDnlfDhTi6Lv+hZX4EnKHEuAmr5
y8yBcJbDKlZOjI/v51P7EhoV5L34HLgYSWLU04DDb1sXpqvTYtmG4br8Omjk/RH6
dyQ0zmTvK9UbdP3Bt7KC5E4tWXkL7qQ2Kf43hT5MjnONMA+YAcK4RVAPqBcoZHJb
G+B0/t9+USIdEX7e821HPl4fghLAKBUmIi6TImUGtiZoybf3Zo3KFuz6DG5LK1MS
L6TsmjBTFKxwpWjfzmEQC7ejiuIzsLhoeZnegstOlim5O08X9Wu/fOotf0iz8QM4
cyw81Yzvi9WP19qfgzkd0p5X6ZBJraIWumTH5XFimRlGL7P1NJaD0+DnmYrWFd0/
PwwuWEi4EVs495T/MuiFV8/QAOXv2nGZGMwBcaKvBoHcReC9ulOhSfFCj7MUpfrm
ABmMT/GD1z95kRdkUKhzUH/rj4dRd+gNaXUK4lWGyQmTllnVOmKyeJopsXhDHk+L
NmM6UKWqkDWgTAwd98UuHE6687sN3PtndlfRTrNCKkuyspjN8tlNOFx1H88KScIV
q91cq8l1/xC8Eo7jKLdjDBA903cQCmwbBfFw4nOgw+eLygH55SL/Uhnc0zgekkln
clNaVmgtvwodjPLXnpP2iEA/pBM65VSg/IEdfCoqcXenBDtDLel4xxq85BfIxuyF
9Ff+2Xk5S7r108tz7uGId/o/ykwQp+e621EYUaftfSdjjoSP/Q9s4rYTq/4VS5ka
4Ej893/m54Q6Pd9ULd3UxkZaJ4nMe/MIw3eqkYYH6zEgsdwp/hpAooJk/OHadaFG
WLTNs/LI/Lyij0uaUUFqqd6H8Yz0jRD4ET53yNl7krkBAxX1CD9SKtNJcc4pGhwo
g33ycfPnThH9ZOKEXtJ3sI4QfLqnOFmN1BH8q5ydjqxXu0LavirI9x31r6VlPc9B
MPsHg/cST+YMGfvDayz36yW0o/LwrMbuhVr0q6kpDL5k0jBguzrswSmjjTE/bbG8
CsSLdZzrvgZj3fOMoFplVA==
`protect END_PROTECTED
