`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qANC8deqgR/mnWxsJ9Fc4M4weVj2EdLIXZIC+lWtRZud6n/UL3Ch/ACAI8MjzE4u
iGK+H/LRWNrQzup552M14HsvYg4blDDpkd2yojvhFHucX1OPj8CtmZFyILCyi2J3
coTHqnUM2atEBNr8Bv1qtAGN3YQngF0thZ+uXi9MvrW72GVyHQrWXvKw/r8bd2Iz
5iVoCZNi+m0IlgqgS5fwZGfQh5RpCq4vJbMUYfgX3T595iJj/5/gKuET6rNoltrJ
WxqnbdRQPtRs3KLFoBHLEfK02ai7TYf8Sqz45dS01mPtphmYtWQSY7Mj1caQKXFB
RJW1pvKBit08kw3rI5PdOXphv+6k/HvxU1zShAUtj7mKS7GvBLpB7PV9ufzLAAAE
wvoUeEN8p/ZKdU4B3Or6kJ5px0nNQfw+nLmRgileaCJIMRKk825D6APsfiB2fZ0s
3ud/4iBk0BsF70Sh0O8h3+KA+cb9+6VDVYwgtb36oI6dx1e/tIdHPV48Gm4MehiI
lkTLwDorFFYjQ9Kt080iuqiLn/qn21IBjBObdJlAgJB6JcHxMjRiNJ8iuJchqONW
Mx8fo5uhT20pS1Ie6wSVbSWPGa07LKko+H+B9cOwYdMwYj3ZvQJmVJUgt62fUPnm
7nNKrnjJFMFhHn2TH4/uTfYjzEjiLiSlITcqJ19eDPiw/mKH0gTdYBhYffpQOAIO
kpBF4plT3nuPSZ2Z32UoFHYy+4CWIooggs+6z2BSkR/uAyhUm1Vy3jdNykb8IVJN
L2EaJFpY83Dy7OuuPKHj1p9x/KSLoTGVVMT7NRgkn94oh3KC9JdvGUJ3AXdrjqqJ
TO8zaFA5m2uQkLq1c18EyRWVsR7c/Tz/3VhT2HdPFkSTyK9OkWcpBQXPvgAn5qB4
Iainz/2cOuw/FA6DZKbx/fPehLllvQw/6Z6JuiUpaoXv1747dpucqvWiUqVIIBi/
eoGp7ucpjRJTF5RFX28XJ5BSjRfW35/BcAHVpt6hCKhrReHUxWdnayLnuUB9ItFG
b/DQBMbPuXdy65y5T/AiL9KOtT+C+cht0rrrSoPaUEg1t2CoEO3FmEJHeKD4Hv6o
ynvSj0erBCwqEjPcxSAl4fIOHTteQtxWyU3ORM1TG6XISHrWdpd8fvo6mzNN2DHg
STHrlakSXUIR/wc8XkIbQzEURfwuzuu0tuL8LlYHYwlD3hK4sn4StoSm6oy6gNMw
eolg2ubpAkmSae6xrn4Y11uOSqlmcaPU+dUQCJZa4KDyqfzr/eb4CgMAEroGSb4A
VNDdHVuuhgo8CbTt53HAKnJg0La7jT44Q5vJK1Dw5OjQU2Nb6dxye8CZ8aHosVcs
6IthZr22uXzUuK29mXezZsdjzmC8seqHV5dAEjV9dz4icjGnNkYvnP5VtzaBHVpE
XSwUWQBady2WrXbMTDe163TnuFyIAqS07h6Fp4kZEZASUJs4fNXABkcwbL41uS9h
MTZZnOvaUbfvyV+IYgDAnAev+WPDtvqfHrlwOcjtTOlTe++d3UNMcIOXfQmBtRje
wyurpMZxGr7Lo1Lz8oGekB8iZdibua1O5hEb2JALT+RCotBW2LPKMdUteWpAq02Q
Gr64a1U4WqmLrW+2H5zhO+WkcYtQ0km2TXJr4Z/FAFjMVvvOq6FnZZzroZzl9qVh
/MYohDCexi/SzZ/pLS7ISahcjckxr1vPEoUFoSwLp9a+xeTZlfu/huP9c817zyy3
NVU/3b63WtlE8IKXCajLQDGZgOV0IKWD+IkK87Mv4mzPCVv5uNuQwIFzUbNYZQej
G1PFzjuK5GlGjhukGpbg5pByXtT8wGLoKG4dmhwkvMMbds588qYYR1ybLNSdc5iK
iagkgdXS7DLJugMczJoAAYV/pk08oYaC5h/Pq0xEcdjVe2j49NHkcG7FjEjvdCAj
OnLO2cfMtumjOXwt02p2UDQC/xhjHq3frXXlyhFNjYYTOYnfzznxSlXHu9WoO1ms
lIXK3aEaqHUQuZ1P5rVHGjVuh9SJnBAi5o0WSC6foohCO6oKv2mspfUyEK6qEraV
`protect END_PROTECTED
