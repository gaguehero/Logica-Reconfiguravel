`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucj5nj0jzEOIiD4TGvXwn7z3ER/yMJ5Qr+IiuDH9hplYC/4BY01rIkVEYEoQSJw3
kXUV6j2oNvF+FJsByI/ogKK4nz26t5NqaROWtM0Dh7X9KToZgFCz3b03B2d9aDtJ
CMZTa5C7pJT8K0/XYa93PJRS8xUHZ2h50qCIycC22EhLNMu4iF1xkjIV5W+iNC/Q
eW14uSR1UVvGxpuL7x+zmSTe7l19Saum+J0CG4ZipRr1Ulwo5m7/hf4ncI2/Ab5W
UYH5FZruwJ5ktlVoOz79x/UkDkCbEGTax9xapoqVZM1PdKVQZM8qz0sQfmicXBxg
V6+wksjnYaIbNbQIL5SL6k2XD6DDXi9oLmcqqdJQnH/xA4Z5nMJ1ktDBfvb+eXy0
nwqpiInYjNyP0ThagCy9IebKEfy1MEnFJvPFr/Px7wEhuzw4Ng/7RB6VzhXoz+6z
JSxfZHI30kqtBY5CO705R2k4gcurt3lO7+beTcNoEl3SXw+GTyxjYnYlG4unOy3M
3RXmqB1907N1qxoIA2gwXdyZvF/sHAcXPhIoL/lmZheVJ9wzWlXQkbfxq9zWTZ5N
f1m4k32LGe1Ce7JsaOEET2lkLZFaXEYw43IEWUvoa8/06UEBKmUWJNtucr3/05o4
fu6eb356CEvmNMuQgvzPDL+0YHB4iR6Un95kzKseb169/afaw0RjGpAeINwGiT/Z
tbnyKjlYUHgcXnerDWpGirROXb3QdQFliDXfQJN0PFFC0+73I17Y+kgU+mivULF+
gC81mZjrK1j4HZdzQJ7octzMRbLPyM5OKEyJDTmDHwP2kgv5E3rdzlj2wBDPuG1q
z68ND88O2QsW4Yor7EIDV8/+abmMWNpGOSlePksT1Td4g4DCiog7K0/OZOE8d+Rk
xDYtotDuGsSKafFJUxeVrQf/EqkBnh/A9ujWXuyKOtST7cQj8xTEdgvxVYOb3RDU
3eec9nsNgmAr4r9RJ+D5uAYBqal7sBOsanA6l2TgWcusdgucTLT3gAdpQHW9GBMl
uslGyMgXtsTqNGu7RIJUm5C8hFQ8hok57Q8yGcEVStf0Pgk/RB6NN0WJ4U2nuULG
a1JApiGITK3wGRCC+NSwby7Pk8NBi1Zef3SSMVUkrdRc6iFykCrCSCx7Xvp4pTwi
PBVNwNrH6zmq2Jh5a8I/kZB1DLljp6VHZn1tqwMk/2B66H5Gomr8ryiS61Xhy/SZ
G9p24aGXogszmFeDgP2Z8MIZjRE+ho/53iP1wnp334xqi/4dltDAE3TR/OY7+b6h
4IHIEOh5MAsGTWb+U0BS1cL4YxwfuGOVQXvJWogySn4XFKVD7PYZYTHCnSqilibn
Yur64JP2bxE74ZwrstVuHQ4wpXnPDww+0MXg+qJXdCRrw9UTb2FFuTJM0BgQ0J0R
35WoKnhM5c7kglk513quRj5G4on/z/WFoRaR/C6BrWqpENwlZXyx9YawsfHFDeun
AQ+Y3JgWUdu9HeuTA1HQRTgRdfRd4D/GGJIAt5fQjtWxYI9QonOxbaoqdFbWzH1V
bF5Np0sqb2FVLt7qAX3WaBnQ8IsrDOt7ebbIGcjjxUvOHJw7tHgjcvbAB9zjT/+f
jiFC9M21ISCQKe6FcsFjAF5EC9ytuX4sKAK8Se3caU3ziuKSfYJwesyh2RpR9zXl
irsgdDGQl8MoMIN4e/X43Gg9K2APOXc97BFpw/iXF6TUTHJHyjzOLDxB9xKU0No5
4ubVWQ8zpGhGN9eX469uANUUxCAbmxSDZ7oIUo7MIQ1rUugZodBK51VB9ef16rKb
BydODWznU/re9te9dREESMAm1U3fnQgnUd2VMoCfzBGtufUtfsItdNi/1L1gWAbA
aC82KkDELJP6z7sMruNpgOLYDd2mX6UnOuITgj+8biBdYl6pbYsOboW5JHH9OArT
QU4bENb4sWzb6CGuAZTVBkh0uNuwpGa1IFE8EgV/WsCubql/NGtgpE8LYbggg/fd
8AIal5zNWr52O5dOXH+VpkXINv1eoe3Fn6QGv4Pxval9HtRlVgRWsreSkpGBoYQw
`protect END_PROTECTED
