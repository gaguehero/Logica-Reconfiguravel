`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gStqVvnnF5D/Rrr1oIZ1l/DhBFInuM5c9sZDVBOqwOl69rC5jWKQ0cyVJvE5XDuI
aB7dai23eH5MVMzBC+iGBVAZE2Md21d5AsWn44aOtT5a/VqhJ66XjRpO8ZsX4NIw
IAsfQB7eEXX+QTzMPqmk80N9DkqDFCoy9SbscdI9FzSiAf7Ap+HhELuXirrzRsE9
NlL7/fdUT4Gr/tQNk3YoXUx1ZmdtBuln0zawTtJemZVTR8vHQQlY8n7rMPV6d+5I
eyQfmZMf4m+5st0HB0UP7e6VjoiRKjda0bPk2GJz8E2TXUhRmMMXtgR6JdkqbC7n
jZr3e/wLSMmojjlWiU0IdMseymlRUO4FGEooFO59LJ8aBaB53rdZywM0o0yepIRW
fWiYlPZeRO84XoUEOs+ROTWpOUJvSLwv7su8/FezUp4q9f903kdPBIW0hvGw8k05
VWmV6LkwY2GGDxkRQsvVMXA6w32cC9IEmPmJzhwTRH0uIVLNmYMtLITrEHqFJ11q
E5H8qfKVRs+Og7IpUrJiDiVPL5t5q+aDT9zMmFtTG2gDAB0QhQywQ/TEtqsnnqdP
YIWqZAEYaRDtpucOAMdG1GuaATvu5ERu1SHOJpDkGIauTjMmO8WfCJdV80Zd6YF6
Hnj/cVcamqEX22mq7UHbGAKeDki1aEdqX5rHSNGW11yXsjEZj7Lxjte7Z34rm9OT
bkHQ3avP4kcXldgBguc7ubE822n8U/kIRNeq+ESoKSfrLF0I1p6zaoA9itHXBFgh
58MDgVlcJRz1eEd/JrpilE7lTuTBzya1aAP/OuH2js8KWKRrlljQRDaFJvZcynIw
HmUEqjuTevJtn8tFSzW+a9sByoqwwQo1ij0KgXpv9xVOUFdB1WTWf0U+PBE53Yn9
ibMT4Yeu6sgC81GiN6hyVQenvLlSGEkcUNQjpHFpMIdzVs9oJaGZmfdNdQPbMAf6
DX3pzF5fqxpZl+GfxBmSHq/X8gM628U7w42bkqRIXpU9PIg5UZ3lRtZIE1NyGMHd
gQO7JLMO3xqnvzrra6vaNfXBqd1Yl+J93EkYih/i5P1B013fYnsLnRUlAl+UkER9
KDSQPG3pBMR09Uk2j+QP57vfyp9WWhCVkLdvezT8tPIr1vSrK3KFlxhfuCrOBCVm
cmPoxExPkyV5mGpr2giNlUQYqPRoSDfgiVhGgh1jscJprBKFzBYGwEq3Pd16Vpbv
JJN2FFxSw9ETQ5t363wvrsOJB/5xzgD0j+jGfXCVffVcwrowX6LKW+POPr77KXxg
cCSKilwmqvp9i54xuUcHfSdJ2TaDxWy7YPq9Sg4DVeZ4VxIslanpoCBsOwo/4HzX
/v1A1EELBf/CmJCT69vuv6GWYJD7ET8flq9j2i3ValtkG07dMP04RytvDzkM6RXp
71SViydLFaZkhQ9tqZoMgRpwBTDH5lv40HGje4h22RdtHqUM5i24lizfsL9bYS61
lScNtY5skEjJCb8jpHKTDhjpUL8OMK8mmt+TS73gAEF5nvYw8p5x+lkwM57Ib/3+
fRxVV7Rtsx5CcdRkLJY98RELS7cr+1fEDUKctcOTZAE/poWHC/5+nGiFDd1DgqDy
2jjufx1Du8jNAtIcKdy19D7B6klAtGUeFYxr4jY62Vae0lWmyiOVPvnaCVvPcQLz
ob9Hb9MEdpmQdKk0hWqwLVrjvAPjJMasoDjX6+AIjc6pIBwM1SHV6m6NGMCeo1Xh
TC2BozocjaI6/cyfHqCEa+JYa8x+/cfkT3Q8DScxxDMX5qxT/O7mmknUBcUBVtLx
RVbP1EHP/6xrNCTq7+dC9X2u9RNqXwis00lko70Dqzt/NmC7RALLYKTirAsG+7Rz
IkRSDXYi5FpRNz5pmOM66r26YgyrskprpiU8H2hnWYDFK+l7BQZYnbrIYOCMi+x3
gzotkScaKIQAmOro68zC9KNhLUviLkSGt50EshV8TrLJ8mlccgnU3ekOoyadNyRL
zBzoHO6C8Snk1cWeYf7Ip8z5L4/S+NDOFySwF09lXsv4PyGMkMzg+fBsDNyyFmY0
ixBOfdo16jtVyJBcmiPQf/vWSA5v6ufWCuNOxoya2szQYsxiurE5Rp1dG+Z70R4v
zMTYW2m4YtjQFXRbiP9pbYw0P6Gy+GS7kE5rVAl0rnfGWFO8hn/28qS8pwaaW8IT
EE3zcaEO2rXT9wL+m/dvY9eaqgDiCovHke13TVVQnla6+QUuBQODVYtZufWaQ6CJ
7yGD5gMzgSqPA1PMknlb3k57LK0uuP/6r67RFpcur4OOwtd7D2DDQZP25V4uwK+B
0FDHrs5ZIF9R4HrlUaL5VIz1tBhf/FbtzrCZX3HECTbAXucLrcPkg8Fv92Vt5+lM
0UNDrn1EN+NADfhLMj6T/MINrvVg2+qj2p8kxLgxER3/5hqmP0ier5iGwOAuFpwN
QDm8AQwh+NsA0NUp3OxOnzqAatHbq+SliYHFfO815OsT2wx/JDyOhrX+a1o7llsR
Cnt1IgmLsg3Xg0TfM5668nat3ideGBjBDzkQF+0PzpgUhv0Glic37BC8VEBc0ZiW
i/5JBBEyg0Ln1WCq5r7EHfbvMXKN5VFjb8rLMT9EivoFGafYdcWJ2CdnRUd5ani0
XgXACCKP6ej8TzHlyht4vWOWh4k91e3b2ZJsgzxpNLNTq420dtrIiLfL/vjyzCbp
u0dUlhORZSk8ikLw+6SgoYgK5RrWM+aUQ07crrnPbyUbr5YqbyEEyk3C53JRi/Db
jEzY05oAwK2OWEg2Y52aY0IC8f0hxBvOyu12ZecYwFJZu3botWj2qD7XoTN/yMK8
+DN0mZJ/SZXYTkD24htHipMolN3w5S50OJqYWLwU+KMixOh53JBeRKW4nsrsQtiE
HJOlfN1uHgkRB9Xis8Pyy4TFMEtHKumsFaDOmxCmRx+jTIzjeuOtJFo+Br0F9VS2
dZsYp0LVfyCktnrDVprg/IL8r5o1H16qSnuonKP5VXKU/8oQQnJ7Vp6GwBWodgee
pFEbFKrjeIqd5HCJp+XUmmQdBP4hBcvSlzbOJMk2Y3QsiEuI1MS9d3Q/KYFbtmDa
FgPIT+abNiTnDD2OILrYwxzdIxVnzDdPkGYSc5m4x62ZGciquk7yQb83EDDFgp6s
mzHHby4u87cPMj3D8ov/66Xecu2oBlYaE4wsgqe69QQH7qM4fGNDDwnSDUQXjUZY
WS6bNsTOrZl2cN3LdNI7yR2+e0vcec9BgV4BmQBAnsQrXxyTsGwHqurt2NP4p+4p
I8HepPykB0cxof13GHriLNUW1vpa/UOQ8U2je+jemcqen41KktMp+QOnJE9waYd9
NxeaC+i3+L8anbjxzC84fZK7rR7zy5MbEbJve6MD1PiLnuKUpI2bqNrLyXgIbp81
xBEXuv8r5zf3xrraryvPN5s+EoGLvTuEZOUWhneRcVIHJm0LYHzzdsQrBLQdQjZh
RRaPh9Y7220VP5nzDv94tyVOYGzF3QoJsTz6+PPiBUPu0v1hZnadsS+hp2x2addb
+wpvsWMmlDP/T9vWkpPLgoGJtDoAVi0RO73+n9EA1h6DgyFHOXtVGmjNrPyXVav3
6suOQyjW4adDHIkeK25gHynAYNwZG0C4Q8vDGLBaD+7TAkEC4ogmAf9KZ7VH5Uom
XEILDURbP+sMz9EUzZDhAQywtwTh2mNfcKoGlymaSGKtnL9/Zhhu/P77xhBOVIkO
HX8N+nuvQkaFYLHf7+a66LKfySOdXGDRE2LsfrFxgz958er8zjXS1oSpNLuZYEf+
GOfJ72fx7QI6KbaUd1aI6CcRfQ48pMS5rXeLVHTqEI4E43iDQ7lh5KI6EG5O24F2
IrX8fM5fcKCmAVQWDmcxYXBSvWnwm7rzbtKTCnQIEH9rG1U7530+RW5FlAr5oCPb
0mFj5EiTSukQj6hu0F3udaZRBYTu+K2PL4weReMUkpRRenCQtVA+jOGzl2noMbiQ
89ITFtItJ2k+4znzwYgL6MsGPPtYEX/sgCwy/+55HxjB32OGVN2kN16wkXJhWG03
idiM8AMybqVC9UOy4bKdby337ZRxDL8i734bUO6eBr1xAa5G8rAMZqHQiGda3JLG
ty5jifEr4JauE3+hxBq0fFF9BYBPqI2MTlc5bM5H7gCF4GI2uAYr9npZiEokEbMl
Xk3KgEDKqv9Kg/RLQuu24nXxFeGmdpYWm/13KB8ncHkQw1b8DrDpZISCHkC3tiI5
L6WPw+UiHbvbWWKv47u/+HbM+rpKt6KINzDSbfIKpEjf9rMdzTAmBFMTUNSuazs4
YbG9cLZ1YSCwCifJ7C7pOE3V8F7qBtfQ86uYlZK4Y+OtfTzVsiJoGdUduyDdLrfk
msGelq6ZSaU5Yc5bshtDnCSA42/BXsC5JCvWjHaPtJY1g122o7ZQSS3sNEnJ7PF5
CNA0JC2onQ52J3mwGzYrVcCMkYDYWKfwxVh+4ovu11oZQJGpNcbxYuyLol4ip5oi
N58GAlLxkstUGVuZ72aYErma5tpqLFv85MLL6VtPccUebKTiYNSfVbOJLnJbRfIg
j/c6sWeBu6DYwhDGbGTQKHYguatObvsVRl+47gXwoYQcvfbubCNYthZMN6m5BSwF
bRA988v2sCsiRu+NrKD9xGkCEtZ8RRTLG+GlKIA8d7aDiyn6D6KCBrnjCoZ/fFn3
I8LENKl/3H3pVUAwunlWHa/aU1+2QQ5eHJanbLc4bR4MUW22gheg0Nh5dP7U+w5m
ICEFwK6G6WTY/GQ/gUKcZW7OWJFuxCvw5+CoTvfuVCwSAfGdeoytQWZAPlLM+Smq
r29zYzK/J2egC1qrIYrTx99SU1PaZFEMwrE5/0c1taiHKibmvrSZaOd7pleU6Jpq
fu0sOQilF/wScZNDvqqUgkf9tBs6Bze0RxuKSGLcj4E1f1s5vnSq6MW+8QiziEYB
DuQ1kacMvoEKP51/dHykh5AnFNbGwgTsQ4F0pSbPb2ijVYgU0U6yijLzlZ8T0Qfm
gzOTVwfC/ozNAXg6PD4IxdwmNy8Up9w3KeNLwHphkeRE2Hc1k6oFeoPNdkX6M/Y0
0ls3i8CEZYTYzyx9jODbNtcBjMsKY7rg1w6B8bQvoe2UI+78UDL8DdEZA2JewEzj
BedWrXG33ni3sbU7of2SjcJ+xA3vawTBq1IS8Obkb6TDEMQZ072Pve6ryGdoaEZa
zT8fC7wP81HuQVn4VaoD3Mmdl5x+ZtK5puzDRgMEa8hq1hdv41tRKmBEfmDcVZq7
t64Dr3WkJx5GU6pM4MLudYI/iUBUJ3V/BNcotFXdXLTJAVN+2lgYE+heofWR4tQP
1do+KJekCednIIrQikZ3NC+q30Syi08JvGtGV76yASuuidWQhcIEVGRf9IrlxQy4
qJlwe3i6IyJxAtS8iLsdPxvH0RxiP2SHaDG/eC9w9EywAZ5pZ8KNB/816RkPpSzJ
ZZXNab//GL8dUKdUuTY1myFJDUmf3AmJZdp4OKZZjIhjaXOjvAF8ILq4imJflBxS
U+mNl4IlN0B+NQLhFAg/LSmDFbXpHAEoRV+w20mbj6r8ZxllvU4JOav1vFmcy0C1
u8j6yRRwOzhb5ChRpZsU3URM+QV9Q43JmJ77OaHMppbve64rc61NtSE6+uZl2JTT
RN4FVb/HWg2qGCu26ld8ocXCZ2EC2KWnlmF1vocLKIM/884Ouyy/LQrb5Cw6BRT/
znVHBgjYUFt6gXFX79bTz7nJG7Qk9GzKB7cURiI1yv5T2Cwo3LMNhJhBEngF2fn8
aK9+PxfsoBrVtJT3J3RxkRNitt6usg+InvXVod5w1LvwY1afFuEXu/nTgJsPMXLw
c1Lj1eLSI//Rhkc6wbRk8elswQI54IDs6f873k5OX96mqh+/nomCRJ2tIY/m/k/l
UGav4/g2VAK0WiEyxojxl2AdiF7OQ6ZD+GnzaoCRNK5Py8h2t8rDlpucoy2lJMAC
XtHY0hpV9DsdKqfoDurMBOn0qKuKqfxshph8VKApKe9rEbu7Zl3Xsl3gIj2CIok+
6WtL6+PfPJ9POOMBKQ9KQhSfWZpJghwqZV9P72i1++w=
`protect END_PROTECTED
