`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7iIoOZ7Ysj3L73KwRU0Z4ItLMdRhJd2hr4HNPJzrT+ZS9cvEgqhZPGkEhJcmjvd
V4fqDfYOna6wOFVqZiY6kI5lg1Dlqb+G+CJS/0MGbEDTv/MriGFjBN1d3zfz70Ba
9L79/eZcdsV0nA29mG7KHXV45SF+H4ys6b3xdmM8QIRiJQWW5TJI1SrW+9zOb7iF
PbRY6jp25CsUPFQzhiAyJAbCNr3HIa5MOkErPHSB9Gq/q9Mv+SqffTU8Y3LgWfFe
cbz0C0s/7EtXc1/WTLElLMKnuQWecBFAdq+dbHmnInWmW2GbM5urmPPRk+jgXsXc
9P+5mbNexzUJ3SLMvhJg+Vvxx7+fGZ46rHCK1DfBts2jX7mFFjwIlmcwcPaMNUux
i6kj7P4A797CY3L3wK3aDDUVHWXpIskctcqVZU3vDg89Fc4NeCxMOTKeBoPyL+0N
AHtavp+I1Er1kFrak8qoRKRGYys5uOeJ9Q6f0Pd5sn2gTGulHcZbJVL/JgkZBJz3
5jTdxOnQhU5+U2Lf3RYmg/HWJqOjcFLnAHNkrQXbZn/O7PItQRIBrCaB2mbV/3Sc
chCrOCSnM2gg/+vkuHQvAi/i55IQUz9zpKVH3x3Oq/b4lZYslECgRBKGw9rwgvM7
p2hCNSswWB+esaNRnJ1D3A==
`protect END_PROTECTED
