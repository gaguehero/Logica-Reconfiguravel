`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R+9fzrrgaaXbzdWBEIlx51rXawVE4M0QKrscsj91XKv6DoT0pWWn52cHzZQPm5GA
8eoH0dEoFZdiVmkMfXWqgmXaD8EqKNYUiPWZaqBtdIXB3Sw+N2nvvk35a0F8/y5H
9f+Y+aerQvsK6JYr2jqzxuKqdSJubWpWYD4uzV6xi/AxbjzgRckcrYytviPvyE8z
0d94ih78HPY0Brs68EIxfi6SjrcghPPV00xB7TRXlPsaB4N2mWZG3hOU/qVnnCYo
Ht8u8GohQJboijoYeLet0MIRrYMIvYjzXU3M3bP/Nwz04RRnuo+aq8yvqAEPPX+T
+3jeTW6whJ7AsbkEx9MN4z6gm4GeVGiyeRe1FytlqETgnw1yrrudDAWfDcjM3E7S
DFeD6lVibKT1VWvmXMqCIOvRzhrA3Cgt9Nt3yEZ1/3bKiMEyqBwWQPDDZCK8aZen
s4uR757zvifm+wUlXol5lu0NkO66aec4WGVNd159NSe1HR7Fb4ySH0zAb1lAR0e0
qhT5Au3aMTuO0ZRIFceJSCIa7IVa/jJ7kQET2aA2o/8K1gKLIHsdc2XQrXIk6oXf
IBj/OluazArwAFRCvaVw74745iAn4QWCXdCJ+zk9eL+qdtLy8YimjEfiMDm/+7W3
4jszMSAwsUi6ylD71SO4Rp8P0mxXWNG3JyD1MkpR9fSUyWn2tQKToVvJPQBg9zga
1CLdwCKgIe8VAM1/QIXzBtVyzi0fW1xbm4V4/mzYjsA=
`protect END_PROTECTED
