`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Suz1Qp9rjXxUYVB5fHRAVxfSkULBq9y6Ms/RRmptGu2XbxUjfzlGsV5ClIfFBS/Y
Xz2VxvKpgNjlRtvez7TlAZ8zIZ7+nkLbQ/0bNDtdSrX/Mroy6tdWRKceEEX1lpro
j6pHKmCOEQThl86rx6qaf8LiTjqT5lOlousqQDQJfql5kW5/0soc5sN6HsPPK29+
k/zuv8ait7OORxzid9PNtemzVz7EFoI8HtP3Pqqcw6fbMfoTo1Lst0CNUeS8QmKb
Ow/c1I44Ey5+/ULaSc+1CeoCa70vqO3eX46fIRpfG449YynxOhbq2b5wcYztqPTX
xhY7o+NsgQhfo6GtfykqgaguHkiXs6eiYXcoy5AqECRZx+R/GYStLb3VsvRMKtiT
zxm4ksxc7Mh/hWXC/z7DOzUiwYuLROizd7Thj9cJwo8orwZLmlYgGsMw3Q87diuf
oi6PDg7iCfTPoF17bGZ3nQFygtG8WkCtq/7EzPbfTR7JOojR7fdoAQYc1srbbuew
8mqyytXAMAbDpwXkl598xxA4ow7Wk/ki1B8Y6/glkXmzP75sJuQW9AZ8Sb5cn0Wu
rZweVffIW0iQZGaOfSPPmJEBm1UtJE6CX4HauidxYrP0KNbr+obACf9hkF46ULuj
52FZiiFjARYsl6XxfY5Xi+qEIF2YpEIaPyfyaGNWkS1uh1v2WRKchJ+NSEbEjMd3
hQHgxox3TjuEfK/coNY6rOT09B0Pxy8ympaHTjz45CCds/5yJ8U5J9b4QbFJm2DO
01YpckY3Vwy4Ma93xkpMhUb6/WrYggMZuHICFETcyhp8NLv+pPPFdjlrkdu/7W6y
nFNc06DOEz0k+vvauJqTbJj2BD8JQbiIibapImShRmwqAneZGmsTa633erSGN0U4
CaSMwB4jSwb0A2uD3LoHEp+5HKZnZ0e+nvM6nr4nYvvISgbcgCqS8f7MMfm2BuGc
sPGIMiWAxRFultttizSv0m4wnKV+O5Zh+XnRpnwyVKhkHJ+u2hMx+xDpQWKewT5l
wqnIp6EIVGtn8WOG75y6ni1OkIMSGVjIkMdAyapKuSPjW8lXm3bdvNvAF+Ep7LZj
HF7nkhosRoWhVwFftk79f14S1B5RaS3tAs+6jVNfO7hunzxk3xT7sHS8KVAfSKVh
Vpt0xU5mjTvkOaWz/RK2O+XH9vshQeA6/GyofgwXLJq0jxDOlV5KvpHDG1zhAkfL
JO0mzBfIzxgGRTZO1PMbvyD2Ueyu1epeJ2CGOiIeBqxFRW8NUVUGOltDIUnVABIf
CedD7KuwQr1uiVM77uxYLsSLQ+M9zOULg0WQBLK1UnYAKOlfxtjeevvtAFQHVWFw
5Z2jUjnkU1DzvypmbKVf5vyo025OjQYpqXMmAU0v+uVTHvIsHfkkG3UNHl4EL7g3
4Hn1vw0d8k0JP067QxeLq5eC4ZHib0Nq80nZAj6/QQ54ObNExSYdIxRsN6/BFXW5
41DxP8kRGmdzM0t8GqPSc/z+C/hlmZJSlBdrvfD+u/pfQUNQUDEbDGI7Wrj2nlJr
FazVO+0mfUYxt4M1fJkQfesK4oiRKrQAvxjxKwCmJdFLAqcaqKyNBBxE6kUb3am+
657TG5Dv/5Tqg7D0tfBx9I28FjlWnpJuDKZtZ80JcdxilPLROd2yEEBb4XyhIv87
gS8m+NmvJt3WORwZnSm8Qn+38/yEoU9/o3Zc5mUD6IgeRfWg/ZFbRlROZLE61OYa
GxTE43jgsJKFxaORlVNdz0TzmiDrM7vRQqLIlpW/9p8my7+jYh0nNcI8ZWRFjZqE
JmRQzEgsJ+VOnHFI8gXvkNluN8A39VFS4nzF9vyomVAKEjNh00mvsAAHYRGuYM5Q
hIRlT5XKxJxqnpRPp3WEIekzenR90W85R2Ci90cWdTa/y0YVRjipgsc5BbOa5z6U
nuDrwYkinVQDoCyQtKbBzEb1MvKI+FOtDUZerdkkiMVFIyxnTGzWfu97YhEJ4zhi
WpH/4uhZd2AUJPcO/QUo1m9RKQXO/AOMDrfcY5lYx2gOwOEmMRfu848vPzTIYDrG
bI/H9QywiCU6Iee+BAnOtUrbvc+zcgIvTUihJ51YNw0CufxajTczmzP1PwcP1dG1
IR+7jvCGsU9FzLFGDH/POAKrOaH03GMcLew9fSe9usaE913qzSA84cDTWZCzWMDG
MbUFP/xTOAOqdynVwuR4mtrpNJiChbLRYHc5RH112Yfz8TovGooShgnC0fem4WHS
AN7mkpCKfOjWX27Lv1PSMPpgNbwBCpLLwHmyveKCPchnZVpL+TvXIS8ajPe/yGR6
1Xq9BFiDljZ9thQUveyhd7JPYh5bsOVybvN9hLvPsFajTOHBEryL7usjCfdNNWZt
PdLj5u6aBC5ZNcedovCGIdiQHrbDPILc4s1qJnuAn/xbMDhimO7JZJmfAkwDwlRL
tmttD0vyKpxRHyrcIWu126ZZdDjUDd64AHH/iyzDfbxl+3t8i6xvMZK1hgi62tUP
J0gMm268SKCl9uYEEHOvOZBpG4+2SuRqGX1yiVfJQY7BgZlfzk+2KVbkej0vtLQm
a6Urzu/HPHynVQSLWujPz6ipKSXbGgebjbYrOpQNVQ3DbmVWblH9OGW/HvyZVstH
HqdzoDDjIoM9MogVrYExbbGZYhOc1Gk0hQJcq8WkVwXS3yir8N4PMkl/aur0hy9G
dT/a5Yta1UNIysMqpfxXn+Vy/i3ycQvFuYJLFaZfCw1sV3E+ibzd9te86d/t6Yk9
lNJZxCqfr3BrCHE9cZEL0qoRr8IH1VlKeKlmT+tbjVT53b+NF6Jhi5k8K1G+HKkh
F8dCrG95DQuqJ1oki20bg1mBl6WI8jkqZgz4qn2B+e4I4BalhxEWkhnwn2tX+r9k
lzwHuHI4pQXd+BTnBI4c+QLMGaXM0T800/AmKLDlU3PHjOa2sUiaaRm0dOhEBlCr
Urm5qK4PYGbI9P+ZpFPSEJEAbkQw1Zlgr0NKZqjoMZpYNku6t4l3eLL8/MKID4rk
wk1gQK5RdH86V92AIh87zDc6kUGW696QKlgTbKG1Ou9Cmh5Ni0QsQlpRzFphKQcb
dgIgXCBDBvXoWuBUysTNdoAwqOkb9gxmGAv5k37E6b3T3XAX6XRRhiumljpqguKV
NjJDB0sfr1ahveGaLdEas1NeEZUXtbpvIxUwB3qI+ZxQlouZfuqtrpNV91o1X7BP
z2gdejLHEgajhWvN498JOdJezH1Wb5HcjVj83fCEcdm4/bGSo6x78G4ECxxDhA+t
MjLJYMtPKndsabPZskCDaHrJx780Rgdpdu3Mx/ZHGC43Dfi6rGNiJS6U9KXcpJ8h
/bbGVDoCOPmGBOrIZETBQ2BignNEuqrZxBNvT4gxnrw2Ewe3iFzRyPKbsB/xGRvw
O2fFWAc0pEfNJy62BcMFrzv5Zi5N4f5mmEfBPSjVkU3v1fqPgZ1DDxiuSR2gLiXc
Mc+RgLOqRI1P9vAuI53SaaexioZ9xOSt1WXaN3EKorlZNBr1crBchaM4JkmC9pkX
B9FX1CvO7Ngj0qKt0FRHJbbKvelgsY+eZCX33xdJNFnZV9K06eYFWHhdITobBM35
HGElqjeavlSy+fbElfOWBr2U/bGM+A2LhSVmjBcJV14CJlmv+ugyA5iAEdf/FQbp
mmyKD7jKZXSoHfdO3Pd4iacr6bS8f/7/t/PAragkbzhicpPwiZw5TGesCzyPA7k/
q+xkb+Y567HlNliYxt1YU+5JNJdR4ajjPyclZo7mTYV1PF792rxg83n8Aw9vW4LQ
7x2iDMGNQLm3G2yG6xVitHvTzP15KfmAg+IP3s7F+5Say6blaN8IrQnNj2OnLC6R
O1LSomLwdHhmjxUBAIPSsCAs6kARgRue5znXHaLHBV4pBfrx2OBlgUhBgIbHkwtU
4qK+TqRYzDp7KfulCJcY0R+8d2tL4zZVYS6e3HYI6HtByq8U0Rw1FFu6tOzslaRv
XeE9wGceMngrDG1pjfH+AvhyE1eSUqVDLeiGzYARFZF5gLQf5Avlc6O9In6WzHbB
2TASjOZOs58cVWh+BMfLDFII7CyySX3vVhYAUloCmzyNZ87G0xpJg/EUESI9yRSQ
moQg1eM1wdHwVJIpAk1q8YpUT3Se/QqURz28tvtYRHRHAIv6SwJv8sj+SLOcuVkW
oKTbFX1tCkPyxa9SsnAWOdf7weEhIP2GYnnkTN9nonwpXRXg7iIXlXj3pcoXVq5n
6TUfk5ho+iZObOGWpucYInlWM68bBidGZmzuxjvt1P9yO/hXqm//4B8VJn+jJHJZ
2xv3aeQ75ffnUWtsK3FAfiTGXM6zBE4Jyw7IwKY4DboeNOTHJWd5o21aBV3nk5gs
ImBVGQ6hmSMMnsMkKng77FVcwZV6I30QWknc2DwtTgE1HHCAT35aiHevopdBgbmr
ns8F14Rkt8BskJdYavpYJUOBKh7DOZOvnPyfVrK0HxnskQ147kCFKhgwBVdM7eRP
GLXfqFUYGNyJp3h3PVVZdTxMF7wNqhB9cIC8WOABg7K+0no5P1jLe5Z/Eq2T1RA1
mPBOzKgO9kd8F1MS+ojl+gBs49GfEqILd5clpDuIGwc1WXDuTNndX1Engal4k5+q
N4RfFFgRjeIbByPBpOc+NlMvgqYI8bdw6VO72qqZ+zH9r2WZ8Ljt7lEKSkNi6y51
q2Rd7/ownEkLFFToLwReel4fVGnkcSur8GVTQ0+KV+oDlLlP9KVBrBTLShAcRfgN
KEwl0esnzqJxm72eM++4AN5c6+RJrTVPmqzypJJOqHc4vlC3tyY/+eeNwOfz5uHs
mUakBw2JDwKBkXA6EtPSvav3Tc8vxLN6IdzpJDjnCkOlU3b7mMCfRg0G+Gp9JAGR
ZDCH7EEAaC7aWm9KADIZEoDEgHm8FZ+7dxTwSTq/LoT2PDPIWHV78cnDEp/tqD/z
xwJfDdHB6n7/91seBjhuba4TI0b/Qh5NREPi3KnltSlRHSwpSOF9XA0wcSenVjvS
+Q4ZvFa6vTRHvJMCegNODKuOBnyGRYy6AilJ6RYHP9PrSP2aEAVbNfuYPjeZsCKS
i04U2sbJ/jG2sTkFQxKBvPRifS/Kj/FLJtBuCmuQ/+iqdDE3Qdx14wjKBoLEJUi/
NOHZkrQaXbPFYDbgx7NDGXa2Ra9ljGrdkowCPKH55z8XrXLR6//zqZ7GN66+NFH5
d6bMnasQ/hJ+srFRgQlo78xUnlt0xnJk6a8M5a1vSYx7tFNq1nS4PMo/dFIDo1GA
h2zimdbfReqCv2QlyCadnCNloV8wLW+y/uOLLbr+qaovdTOFXBlnX3+n/akAhaaK
alftvbJHUDklrZpUn9dld3m7oYbV2OZ2gDdbnj1yzy/gO1B7FwS7FrgDrP1ToDJt
QgFWA6pQ2u7b0qomUzHIVmNHxMZrSbn5Dpu5Y11c4Ulvv85lrCgelV3bQ6Ect4yN
tY7f34sEsg0mduq6WPZV5SOnNASY47KCgb9k/wJPhjy000iucsjqCfApr59rKIGX
nGY8uDlyd9rn95HOSBRjjhsUtFLSJ8VP4uj+WaoKscOrza9uW4/T47tMLuwh9is8
GDVEye92CHZx91aaxwTNVjLdStTna7DGvSurtldhc5xj2KIaqZc3I45nsOei1G3S
w04RVACaMog2DZlijt0k+zdhFshqGCrVxD/wU5HOgpkdSjknLZbawexO81W/zFSs
mt3VmXaUEkpSMUnuN1UqFNwG8d732s5cikyktCDwniirdBt9Cix19/nYP7gwkWLB
jcy+AUNSMeUgIF0ABAJ13Lg8NwqVKVbV3Ub5NrkiJpkw/UU/DNygIOQQ7xwBHXQ+
OnJrJ4vapNEL+4oYRXcyziCNJFUn6E2Dm7hPlipjaNg9sqLvgdcPRwHmpGOvLmI6
Bo1IOZot8USO+YE1PfqNOIUFracQAUo06kgSpmM0qDpRs4amLiVjx5KVwdZDUBbv
+uVkQ17NLLWFDnjlHxhXJZnQt0mRlHdLmXhCd6A2NQ5x+HcvsCXpN3qMEK/3IIE/
Dx2y9K4ilv2+XHVJ/gZi6/mrHHDSqcPV9te9ruSSJApKTAf/eVM2M7BWp/AGdzZO
E7U8bwp1AaJzit6UO9k4RIBjiYFd6/JbSx87Q6D3o6OCVB6utZ0io0NhMvhYwItG
MGeeMF7PbY60lIpg6zLlho5a9EK9DTG+XQdLAP/wTBOcrW85UirIBht/ttFRGl9I
V42i2ofT3d7QoVTZcrXEe7n6dVyP2XP5y0OvnHbJ6u02VgERWEvnIDJZVLog5nvR
umqejSlIpYmvouhSIAJWEDId2KfbPhRu76tquE25wfOpVe3vDl/xG1tSKfOfvERW
kV1kPTzVErSpVPOQmQ0YLYKtdd8HAJzuUrq4heXF2cQlqvGnFejNp0HupA04HTqk
1x1OfwD4OgaC9mh7pq2aKn4Dau2aw975VBL47Xp1AYH0JMzE1BBDw+WExHSe/EDs
pb2+G1lIM5DoYXQo4HJjI71pclGFcdVVKQa8iJwJf6N69vG6+C8874ibiVv+7bCY
CCuu3Jk0pExXgt3mhIG+yIaBfpbBgco1XyFOPxHBzCGUTRrfi7bzEDvLJGxxVutp
FqPiNwRvIfhseyuepafHxo1YUV/AYSCDAjLMhdlDQbuL6SdReUo3gsapEUaU/odN
Yh32CtUXkZpi0p1qAjxEuI2DrgCXqVXDYVwY9HmfuSwwyayOn2aQMeiI0hMCkNbA
mxBg3bW4otbDKYcj0jkGwVzu9JhdeoG+or5nn8uEfuzu5flzof6/tcY2avv3R3cq
AKiuWHO/Fo0zz4Gkh/TMN9CQYAFQBDaMCNvKY3KxFM4MYIAlkNN80kNuzaqnm9N/
v4rTJ5mYzHKjDtLAqLverXmASBrxiNNAqJIQexbd09hAWpm4DYpIJNLONEPtsx3z
q6sU4437frxoWxD73oUg1mlkj1bh0OMWpiBCg2bsTyvkqoBiwfoGtSY0kkyd6xgV
a2FOfDrzaD8JwZ7X/xrAAO/S/MEapXJvrzhcCI1Se4+AduZhWVgWRE/tRtuth/WA
TSlYWxT3si8YPJ0IEnbhLLzKh8I9Qobjz27bfkhUi7ZS1iroKRsBUk4yMnkumJeG
QqmFwV3BxunkEU99jJQHA4H9N3Iycaz5UyucMH4PnbRy7XC5BOWMI4tgKxZ5t3Da
Jymxkecz7MC9YMuXGkBvN1aGqV8VmY+M4EYGik7QcKzk/MWZUtbm+hhmbjG4LvCg
K+ez592m1snBWW606NLvg+rfSVmodO0iWbX62cGREf76sFm25lm7n/+c/RWDnaft
StgoyKpSvc3fBgEZwL179onTTjN81bTzFOtsl2DyUu4Bnb7vlorTKXwdAR1AwN9r
d8dPlhIrgM1/5yCxMVfQrI2GoqC2iOcJeypLBHMRHcPgOZ3ZWImnXa6HNftw2631
Vnr1v88o40Idv90lN8NroJMzeB8PRz+DaSjewSUzWa1+3jci02k2Du+AGjiCeawe
pMq43wuuAa3B8EedDi0SKy+9Sis1nKIzQUmQdWKCZVB9NpVM5B+0gsLGJVcpSGAP
ZG/tycfEpn0tZJfrzpaxu4pR1Sv/mPdC2EPNSNNwP9tvpHWXx0s56BCUaqIcdcmI
9L/uxNFvnt8dLnHZDwlj04sIBWleh9FY2jX1F1BlRn2a0j7AIH+GWWDu/aZYBLJl
`protect END_PROTECTED
