`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9V5eFpdRnBeu/7k/ceSDd4Xlqb+0GtCzMixyQ4PtYG/ERad7+BstCKO2IwTpuHzS
B8P+69oSrgaIszgLpNSyqA25hzxWf0zuYTiOOz+jZJofKrPEQ1REo68quzZZtG8w
d9Z00aFosvpMfJ1oMKtXupyTfdQvDoXp1wsT2ZOIuCqxUqxPRkdv+RkENv9xkXAR
9oul0xs9KB6mq+g36TqLL+/8OKG8ntm23FycngnfBPUHBWadf96abl3x95h0BhaJ
6UFnWWEeaZVO4RIlTKHeQSJVCXUdzguRF7GdssU5+kJjkLk3E6KT34TrWRNjlDKF
CvikVM052i06g+GIySnndeKjhg6KbNziyJ6VNz+AVsMAYe+3vpPfgU3GHgyhYu7n
0IRpJjzs3q5LRmIXc2vWu6yB/cpNI8LpNlJSev13B+B7Df8hqPwhuaJTNHqSb8HR
p9ISyyk9zl8/sgqxBJcmZQ9l06uASKqRhVemynY4XPEOouiJaVE5FAPyyt0TpW/G
qCQDdQKHVkhFbX8RKEg0qLBeog5vv9ZG6mkwjKFgd1iO+bWFbZkbjnFEPTLyLJNB
ek14dNdFAHYCH5GLIV+3a+R85dNlM/VZtC/TCBuxzlDI/b7N+Wki3esJXRnmMvX9
GZmCRNxBnCNc0RVRrjoQO5I0oMfUp7FWJAQXfY8tNkeLGOmNs3d8U69cEkc3Z2RG
A9Pyf7jrexfPBwp/WB6DvkmmKK8smxR4iHHtlEwZeH2C3CWiwEnueeOCXhMD5fc/
mwgTsoALL0pF7hoSVzch1hkICO1ycWEsQG1q1YNSQ22zNCWzwtIBcGZObGKvgiez
RFubqOnka5LNVUuq+b6awvCFhSpknEuuUPXEaYZfgnYaUT1D8mevCZgwFfpXea7o
+b22+4CRhxMW3yhemwl2EdFz/XxELsyPo7gMaiYEKqvkcdp+S9e7kdw7TdmRU8LJ
cwxkgv3PDksObUfdpjsE9sckROLVXv8pIF4rnwd1L8g6S2l1/gMgGuQNXl8QCFNy
MSy9Puh2yv+OqVt/lpvz+oirBBjBkXF0Uw1hB2zcRZ525pyTe94tLdV5RZz3hcOm
22byDN6Zz+lTOxrZpXPzaAwaz3HoJJx7+GQLW/N/suKN8+MMkgPLqiSQ1lXLzGgy
1fnKKYLbaWBphSnZ+BIxfYDSc2Km3wirAny81hsU6eATlXgmhhf+2ENSIpXGl7Me
d+JD+RJBRnYx3MvbV5UF3wsU7q2pBmPcgPlr9vymIRiK73+2iEj3wJOWpdEfBGR3
yj4DD9LhVlIAUpgIDlN5G2JzMVONpRKDZ88xMTcMNlZdonhwEf3xSvzdsHgN7OOS
9wxY59RRLcJaZWS5JruhWx5sH2CIPSgNs7tnTlsXII/lNwwDLtr+6d8FJ9Ip3mZG
oUwZZ/KiyF5NpXkOdRvxO+utlDjs5MT7SjG5D6tiGHkYXSuyPiR8Ygsrx2mIK9g/
b47tkizEC9BIzHkI6uVzXZglGVoL4hGh31u9ShYBIdctdeOCay1Rv+i/qIqQYiT1
tFQCQTnNguqp1ts4duwomm5IsKUYt7mKBoIlPxRTNg+TwhC7+7ZMSeM/Y4kCFLpc
SBepdgKoTSuaM7QWuxhP/8fZusu6/fnJ3Jd6EPOl/M/NTmdMNdpSLT1Ift5S2l9l
71kOO3QBMQyYYAP4aQufLsiWpXWvuO3+fJrBaWOrEuXUrCj117rP/9BIDwOkl0La
yh4jtw6JVdnsaZ0NMvRUn85eZWcgmLl56gZBeUWmXlxJe5DiMpNjG4ScC4Bjdwdr
DYC6tkWQdK6Ts5vL98lUXQ8Wqf5ShY5LBikFC5ZRdQw8cS39w0WjITF4yVoulOps
bKPu5GJ8/YPgMbpT2vSf2l5Z+p9Q2Tub25YOi69yqIBUC1paaQ4hyJrucRM9fWOR
IUp8mxlF1LumONBooMXUkgaypBFCO0RGpLGGU18gl11GiW8HsybBxxbqts6Pr2cQ
vTCtAg7cLlU6zAqoZ3rRROWZOCIod+CJDAktdWSMor+snQHo3RFvdDgxKpYijjqx
sN3GMWAtwbXTe8gddC2fT1IBkbtOSlamoUpLpOF4dPDXP75EGMipZwjWq9YnP+ZF
kntRkvBz65zgzxi4Ne/Mw+kvk3kDt1FoJmj2ab3Xj5SPYqy71ZwFwCK+fcFrXQAh
kTtXYIoMuiDInDQPYTTNv/LkKr6RxYrGEcD540Y44o+G7KBQMPkjMmYbyRAZw68v
eXbGvnxaMrLt+7spnGH0uVZv12l11N/iCGwZnGxq26wtdHK/FK/AYuAHeNlu6aSI
36TNsqIn7LPIVdXswjFs5wIGYaxODSL/zSHi4cmBB9QV8qmoaXHgODRI/LzwhoFy
COlHcaPu++sJF1uwkVXpYFRIfkR/Fqsgk5AxmhXEbncVSZ84ud59RNQ8GNQbwWOh
D2BLOGr4WAET1inV2JR54/57FpAKBfEBamS2eP5q4j28IyQOmBQZYbsBK51HJ5Zh
GW+GCIaDrj3X/xgO10uTrURLaV8WlFGWpz1ftRCDfrwByYLE6koSFY2rX7gPYPH+
GUX6ril9gUo4pIKbOQPXMQl8yIkY6XQXH1TE/+LYPPp2RunHn4swge53iIzWEYmR
eYNFW1AegNNTXMlC4YLnZx4pTB9YXcxKCSNfA9pO/QIPqaKjVV2/WfpBSXM8AysJ
hNydjqbILhqhw4D1YrF8aItPSxCk2m6RCc9oYbY1uHN6loSv6d55Gsl4gz2RTYMp
iQzhhdXeY+p2bUO2U1Y12S0cKHCCyM8tEUFUgFEZo9gcJxdQY3Rrac8lD6LfT44E
M/acQppDUMp1riB0aiMMyAdKVdtwBtBT51rcUA3n4WWFeOoFnFj2kxSXODLZF+IA
Z/hjlkCKYMpIHDiwrb+0Z+ie9ZeD6s+PX1eoqfI5CpsLEm9wti2MebjtCvWaugsl
5Skic0sBI+nCZKF9Lciqav23duVzMW6jSAYWxoifwVRgb+I0I69JM0lN79wfQMb8
Pcp8wf0NVEb6DnjB5O+3vi4BURGBirPYbw2xmtqjPs3Svol5LU6qJ3IGYMEw514x
iwt7XfoLwv57jj8YLvlugdRUeWShp2hFUmeD2Mr4tvk+k7l8h7ilhZoSIwvSv8ea
os689sNeGwotSszfZ1j/ZN9Ih9qMlVYGGxvmGfbGKkhvHIluftEq5h6NbXrlUNII
5G4PS7Q6164/82eQlaZ0uDTsMCYA4mA31Zson1oLl4+j05GLg+33M6NBw/destaH
1yeTqConAJ+HakSPoEc1bMIJbs+woSwz6AADdX0vQBdkN8jVsHOFuw3dcVJay/Uj
uy1+dH4k43rO2rCI7NBqwtMDhEKkMl9JDfBXYdlEnF9finy5RmhAn1iO9xpGnP7Q
XVuT5IEDL6T8pOrUbTAL/nQxYCHJPWKJlin46SefXN0j95rZWKjUFYLbQuRsdbLJ
g03g3OKwWGgvqjY+i6yK60oTsO3SLF39/XAFxiq4cm7BnwI7+jQZph9bZJfVW502
Oh8Z0M9q0RP4pW9THY8LC1CQ104yNWgLmSFsd91LazeADJ/I/4UEx7eXmkUhSB4R
m/70NCMcKLQ8/0HczWUCHFi0IiOf7pyo1sifqOc2Uef6dwLkLEdGKZ+Ppj7KekSP
lyMz2TJOrYakGw8wsXhbENcG2qvimhmEJUgWU3jkcH+koS4G7PFb7YbpRAVfwH+M
Stgt+dlWZgnlfyz5YyYAYExsozrlTM4mqKUy9zASvr/q5wr71ohrAkPnIJXhkb0p
6OmKFAiE4Dbk6GNa8ICbUb6k7dQSexwIb3rngAcLGuckriwO2vbJCRvcr/QtkVcV
sj6/xaYkDHDPrbeW4aNA2TpUV+/NtRilEu0aj5/xqj07ZsXquwM9FVQr8wxdBgEb
6haMFrgHc+2fiiVmlomkn5XafCO0lTw1rQZDLc0Bo06kfxrfr0n3JVrSG9SoZ1vA
i8+gr87w7ec6RnpUmlUqvwvPbZbbzMWhIAU87qDQeRCxEAkoy9L5kyWrAW9SgQMy
DHLhfSPe/w9O8OcahYyza3omyVQ/Xj6ytIIe9KXKcKw+U4aJxSVFDf3Zgk8223BV
PEduSonAyeubOlsPpjdoMuwM6W3HLZyS5UF2tzJQMFSPXQyPlQLQxRfXv1f5WePI
e8DjfG9r2wuRVNVgntE7H4POn4szmRXPrSxPa6CvgLKgpBbUiI66gVd2PEUvLUQK
04pmUSDZtU4ODvpTiTQ/URYb7n2KOUsUOUlJ7dAoGHfonZpOdGbY2vClcGC6Jtzk
iftlx964aqN5W9O32lWj4+Abgp1QX3JNm/jPhZjRZhTaJJnQNYxK9J/ay8e9+NGB
OCK8Vq8OY/wl9DeRA1IVqd2VBJ+JzqvMdw7ucYCFZdzqnzjfknUjpmMgbExdG+gJ
unt+NOo5xVIAEtkCcLATfyi4hzadXGBLYKlzocxOGUJtsa2EI9uZkWrErT5IZO9r
vPTL8ARD12ONXjXgytkVN0UEPCZCQl+hwedx+Wy+VB0FQ5UYs12cJe5nbm6CWJx3
i7lE0nxu1zggEvl43WQMAsBKoYXXRwmfEyGhV9qV8Y/xTAnlPS8+caLLV1xUwFog
RsQi28yxPvgMcrxTs7mn7OSu9pIY0q/6ac7WKCC20a1DM9vNm0bY7tZ+6yNocOY0
42Kdbt7WbykqitdQMsF64lTgNnKpnTqsPTc+ym6RXqUz+A0v8NIwUek/PSl10X2N
O69y/AdTFZdM/FY2Nqy/J+LwdRdaLb2Bb8EKcjHfGQzW+hBbvFBQG6WxVjAmWrTp
xU8oY8T9yl3Sr0jLqKp+cLS9Wou7j7H9w/idSOB0V5glzKKRpuj127lGm9BClIMZ
LSiaTj8utpownonACMEOSezNff7x3SwfLDjG/GnVsYHKLbl1PE4E3p+ei/zOy9E8
H5HGkl32Tygu1cCUr2exzNJWoKWObVCxq2HD/dOk15PLtDvSVHIJHNEjL3FFd2rP
b1tg1F7ZS5s3Qw0NLVQ3D9TYN89RqDAKSP4fjsiCEP935XpC5OX+RwCFPVP1RzvD
hMpLoYLxJgtI5trBrKM4SmZGsMVuMvLen+z3rwddlij7iWzyvSpyLBXEQVanIqSU
QlxrpYsFCObB16treCrRuYVgfFMuxaNj7UrpBYxD4Gg/TXsV7M90CPzCT5JVTntC
vYYolAc0nxnKYOQAKotmaGdnUDbihl19AE6PXY1+Nwn2iTmA6lm6Nwgx5M2KZ4hr
ChxskShfSIcoD37F+prb7NvK0FoehcNVrns/FxHDTc6oaE7iYG0zRBiSypNR8xov
qkokYnC7pO5ml3vSLYtHmKXBOy+rcupXZIZHqPXfF8FbsDhXmlfQ9SJW89WZ+WaD
tVR4ro6Zvqn76j3qcBJ6dfD69mu4yQj0jG2LTlLDJTyVXd4seJGJvy0iaSwGvE0u
yLZZjtzh5er67cVNwdQMB3uQH0e3xx3cB7DV0HeW1kP7gtnkHBn+hgWAs/NQAqwc
ZL8zY58bAw6ZW/CzsOzcOXHoZpZn1+HJ/Z+9C1cc7YiwatnACt2Yb/xnD0ZV+koJ
6FlHBoo5/tamID7u5jNjQUZmI7Bf8tZmj0EME/4pJmoJtW14IIR0iE4aD+Ncekjl
9/J8UCwcwQWZU2AjQMVthMgqSQDhFZujfK2dY5f8biMNEPRyqq/C1uNPY4SHSHWR
kktC+gPgTBJWEaESFmkfDQFx0qVuDoE/dQmeR0CDeo/Ro8Nq7UFDoUeramF7chxd
nLqyc/mc6U7VKJfXC70vtY0w8zeM1oV5lTeXkN/nEhunbfYTF9iVNbFeOm629gyy
qBkp6BrpEm73OFwsaIAlDZzfQzi8PMwF/XUJz+BTBJwhLgXgepwog4rQIqmr3ylS
Xa0MkJesoytZqgOxfpag9uq7M6GvwFlhXYALeXp1XMeJZBRKOkd2/jrAkfYJEJv1
6eF51xFBdbeD9ces+NebEJUqBvORuftYgCQaa/IniTTGrPfeEIK7rPJXgD4SN4/t
G8a9BvGAHTsrE9wwalm88Ls7vbIxAMfhIqAMIt7906ASCFbDbs+vmbl0H9R1WbMr
5kwZxCbSr2b3zt7eryl9c6WE+MxP7IK79/s8h3vK6kVyBraElLKji2s8nePgpshq
OeQbCDGTTyNel6oujtJ1QsAmDUCCTdoSUQ5RnI20yh51qpoAD6pmimHNQ3F4nHeW
ZLpPM/McCcsa5Nejv81JlWDK0B882NC7kT2DbXIU4KbSezYy59zlrCkbMM/VhAFR
Wt1XO6Cti3CJ3QshC/P25nDzsVEmpev43q7AumVulFopH57kI8+VUhx8X5KlLCnY
1V72EQ177tFR9bo76VWcSyp5SDtIMNLHfanFTMWCAJb42/8VD56Ca2iW0dyIHCIB
rTvBmL8qIRJ+qJrq64H3ZBibosevDCDGKTN9NuFcfjo5mSnweiGx++cshrJECj8p
m3hH0y/lIp7+Exqq/v/ml6Jvb5eM1ikZAPkwTwX+ZXYvO85eMSK2wOg0y/JXjueC
dMWKdgsaC5Btr1ADrR3TXQlhh5Ql53zEY0zMeiNbgSYxXOR/aGyyjlDqFyG2KEwX
sR8K9y9ZB1xInISCgwhffG1IZzTWW0ROlB8DmghggcdASe9NisIr7t6tEOg2wsdP
RZuWwFmxpaHkOE65rqLb4o+P8URbDy4RXpJS9+zfJRY=
`protect END_PROTECTED
