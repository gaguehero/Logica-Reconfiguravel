`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2wfYIk79LoGZUJfpzRQgWXWmMLJ/4ItjCqRGD7fu03oyhnCVNMH7lOpX7hK7N7ZZ
aozdx6m5eWxtFlscQl+Uaj4go1Vzc37UXls5m/FZlqyuniIMWX2dp3rm9bCRZ8l7
h9IKlWKA/iit0KlCBzxumFqYsJbnPPXaLwqSJPabrr/KQPlOLYfybW2D+MWxyAuh
UtToiCrKHjdNiK1VT3pgiHWYujIPNXWav6zyVeeSKeIoyKyzahido0VF2vwU0MO7
72zFW51mMIeOG+/47k89j4FEFXHW6i3U9PHrCxarURrPVHiyGg4Pse+6pLWA8Dif
cpIE8E6ClDOBw1GXQ6O4k77WsFOVUtm3KuqPZxJrno51igQ1yY05Mkz6LCTQkCP6
5FZ2yTswncGQF2i0eqjda1phYcwg5/5Kr4Ipfg0wPEjXOC/XZrThysp+D3No4U6w
EfRb+qWv8M9cLC1kTfRiMjC+LBn8iOAXLB+nVI2L436OGkzM755/9S2TuqOjK/rN
VRKgVcHgh5jlw2pOyVSyFS4GRKc4OSzD7atz6PUTjG8Nqfc4X8/tWbURrlk9g+jy
FLGCtz9IQEYlVJdBYXA8X+TqHZ5KbTAyNWLD2RIPihwCgMta3Di8CiIpe2+tlV8T
S5+D2r+whgpGXZOZzDg4IgM4rPWKueVO80CfsO6jyVxWttJoxcloXC+qQfpCA7fz
s+jlrf4xWoSuOfII57haTlAos5MaStAoMeE5I9tD+RVFD9+AXWfqmzGM9MEb/fof
iWP4VBAbDeIyJzfX6XxcQYv5zNgeGHSFjqld4/jmReq37ZOVtqMyhM5ekkzRO1RZ
1gAhlO5JHQ73+11/pLHiL88+4oW7x4jpkPFqB/6Z7fTYSMh+0E286MJ0ijQy5+oR
iMESdKAA378kucb7xjI8w62v+1FpLFnlz0XD5I1gxQy4P7QFYXNNJO7Ue0kZyGkK
/Xsnwlw9g5WANLWkzumOyoHspaYSQQwxyAAD5q+7yQi2TIT4CrgbYra/2Ns3Syol
iIUflUL47uR/uFWnHX3/wEKWX+G9LaxyNKmCApvGzVnC6jN5skNSkLgxhH6I7Ck8
PcqSWvkFxfVm4JV5N2qZhnmdR4Tcfd5Cj07Fs2O744edtx76RItUUV04Be5V3c3b
fkLCVuHK55l79eaaZT4AIyD1PcYhiN25pXJ1KvOvlxnm6o9t3l4iJDM/p/h99xz8
f9PbAP/2tzp0cKsk/uR6fKT11cDNxDoYZ1e9fQqsBPW5+ueyzncFiwXJGKMCbAz/
sK6PRSDuGPxRm6bG3n3HWQdshiR4AeD4xzFV6GMJm/6Cc7uvl5Klva8F/ckX7t2N
euNsBdXD5tpA0ciXJAv1ORrMQmHipqVuzHCVO1TU8G5WCqf5sSNkF5iAuWsxpQdM
sDEOOpjWPR2SO+9xwgaqMIglHZrHhS4p/2NypGHVgx/mffWs77tjYwNrpLwZhVOV
NlAOGe9xgzHr3NNxnXgr02PBrMEARYonEr9WiS0uhYVxLiizDHNsbXsxfDC0tLiI
2yo5z0pYjt2JxvJSiSMuEXK1wKHXdyoCEcu4smld3BlQtD0HRCZbKh13kPWxyIee
qekajDeV1YZfi3Rx+rgwR4vTwNZ4n/Ormeh23nwRdGOUA0hzJvjoOumWsuVW3e74
A/be+LrvXklEVr58IBkr7PF9GdC4TpuiNLFhOKl9YxQHE2eJBCHrLfAYfDjVjI3A
ojhCJQ40ommRaFpYeZUAsk5gQMmJ8Jac06KRBO08RM3qTD0yTLXAv5n4UvgEFEWW
32LYG5gJs+iSj46HIktlbN2oaA1H0zc+rnRLpgcsRDgU9uIa51VVp5vVhnUAj6Go
Q2X3GA6nNE1xex2a6YL2QfUivakXz37F/x8uVzAmIn2YTKi1oT9kKsRRj9fJtlnM
zYiqhIz+McQgowl/wx3MrEwM/dv9+/XlWF7/HZzY5n6p4+e3+gpviqWcjyMnqVPA
OKbBcMNPbbk0RK+I8ujKdfBFiOeKqDICtkH2yJULZuuuvHdEwD+y54fjHkjSzwyk
ofi+L4TtEpH99IoX1pQlQPVGvsibLl1xboFj0OQ1z+mHRSB8/E1DJhYvyi/N0LXW
yEQ1x4jlEqiln69So9LQs5HcdX2Ungjz6k4mfc6IAhLATP/m+a98ALDkFxKdgXri
Qp1XmRpjyaLNFnzZfx0VXgxIUq6FU//hfnihCSpHDjDoMiA7hwrPNL0x8XJtVMKc
9q5cN/dKKOOF+SHIbTZXaA==
`protect END_PROTECTED
