`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8BAvDsMv09IUjFlxb/ydezn285DJ2UYnU/7Nt9a0NwgdAA/TE3iAHiMERKrm9ir
1bq8Wm9qY1LO09dfMogXdPu+xkF1Cz3fqx9JImQt/0tzNT7EM5f1eP3gEDVVzoEs
JYIF/yUygKO09t7FIejHn/MLMDGOEUS9x/UlmOOgbsiG8LKMWQb52YHZZ5SmCGMJ
LXq3zj04sPOBxEBzP+ZhlamDMIakrWUVvs6KXFqjLHqpTwL7DGBf5asIJzwkTv9E
OYjZ3KgpaS7TsZMFewotxJdd+DNu+TAdXHWx+ZmqcYYVGOBJ0wMOg507V+RV2YT4
ZMZcfUzUY4ELA2Re31yEA7maF8i9u5B/h4sMf3SIbzXAhLgVPxuzr+gRJZMu1x8e
nqKK/vmscbH0UN+s6gvlbFr9Xt8faheZJXE02Ezz8wvvpwNUwv3t4Z/WcKuRAmh8
I+SqQdHpZkCixINyNHT8Ov+ZAg36uCmcULCtOo1t9ll1nn8c2xf7PSQzI4F72iSp
lr+DyxrHIUhSHCsEK12CStKj/5Ndk4xtZEVjG4BFE7L+iyb9r8I4k09JftCJ7DIs
Br/l0GIGexJnFIPd8+38DQbI7qVm7ZpqvgGigzGoxZyREqqf1Y2MpvReqa4VUIIR
eb6nWHg5djbBEoyR/ZB8MuhNmhGOlJ8fhg+k6HdmNR2dFmVm4agsYZ2gLY+4eA8b
invGTxgp1C9JJ9+b57VhuJnC68v91qWhV0CNq3OK3ss9kg2cHVIp8pUoKP48gCxn
MO0frVP9d2D4XcmUZVYxRZqo1LAXadu6yZZo3+5LSkmJqpLO2o7eAPruGGAReIIm
E+TSvDSQuLDA60ZX3fxWqdMXDBLNyLnbfo1vUzVyA810MXu6Tgzb/uS42XxiDShS
alBBbNkeJ6EO27Ikt1O472B/RdeMYVuMtm0QO/tZQ0ZYJTyDD6IvSO5FzjYALEkq
A905pjz5sbWHLUhZ8wuEJsNAQyYSD/cAwTwq5V3MzEybch/0+j8HhIBjDuOtOfzz
C2zXe0gyvqpGKKGY+YZX0BvYoFndbFrd2rBKqsgNuH4G8Lt8T2iHeQOZa5YOl+gN
GTdgTixbm/eo9aDDuhud7dST+rDwuR6uoyksSmYGBpzFtXi3Rmcl8tgz3x3kuL9D
qMG3FdLjh4+8sDHC0JnK4ubHDPnuP0z/StZ6xBbaKWbCiVOaZ9gGZyUqTYjCbeWE
jQsJd1nSYL9Jc4Qva2AXgu3vyRWu9BqBpwlP4ocXRJjDl87qOSd/FpprVxoJYUbJ
uMEo0jlX08pQ59IsTdTRCvZ6PI1SZKmwk2WjjQXb26AbEL7W9JHlJuJrfytmDN1b
iWucbriVXo2zV5O5VoorOfGrNTYbLtUteHxfG6lzURtcqg1F1WDc5KJzdXOc+VRY
eaGYbtxhVFe9UtjJa+1T5RkIxYa0BnzwR4DUsHDgCNGX7okvsAxUqsT3TpOibFBS
F8n4e9/R9i2hes5yKwWICHVq7jqlx30jWbbwNfDqIYuMTZ645KIXAV18cKerr+2E
3KxJtjjEXSRHaw6aOtO2iwCzSDOZsZOQ9kRG603ZmPREdkIezFdH87iK6Z6YC12V
xhBQq3y2Nu6pR1x8Mqi2zYTJImSMzR+OpDJqYgwFtzjK6KHPpRAhbj/6QSNsTae0
90lbqxH9iZrkbbdyRBdLZx8uAOOk5lkWaVO66TtwSC8T9DTsdfa1HB6KDH2fBrj+
a4liyyzsYCcrCKb0LSDbYjEbtGstQ40lDE089rr17jQclkXsHC+Rkjwj6HXwGHNk
JZzdAtAzCYOpMcYcynlvCFaepZLTEIxyRLwfy4WRpEbOPAEZnFCCkOA0kOBQtzbI
SDiMGlwqiwcq4SzhVFBt3v0dLRorMDZhEM5YU9QolI6kQoMPxQRjziXjnl1vZWT3
O0PC1XHwQz9QqR4HHEyjTZaxM/LPxND2pmFGbKW5WMyeEyLjP5u6sn1fBLtuOU1J
Yj8+5qv69K6F/s9ffT3Hhw==
`protect END_PROTECTED
