`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HwwdAdn7W8/WPpdphu59FZIJDesbcNg+pTcjDsICh4NYKw5BVSf4EeiJTjTY2Hkr
c0tQp0vr5fBgTgk6Wh1mRsq7Vilw5QLmtZx/UWJBG/aE8JZ2MRuC3qF63ZnCVOdM
kYLGCgdVtHEcxogT1dB4c6CLr0UnytHKy5DuTklgbaTzZFANdLtJxOjC1jfOmCeH
ehRHntX6ydMsmczInAdYOmk6WcD1p1amqXda6dOOMFWA4xwkVSF5mMJqCwU819yp
4/Np4CORYov3ehftx9jqj99/V/vlpCxverQ/8g8gypKPZk3hTuxAe/T7BzS5GxIi
kJVi5+IAHvx+EcpckxxQLzhuqiY9DXabtGVb+N65jfVV2T+dCyHmdq8OxB/WEw69
+VkO3KI1nwVaahP3TGA1WShMNma+AkVEpLiBLeeYPhoq2A4ibWM+ZhFDpPETfwH9
FV+n2Rg5luJOqxn2dJUKOHdPLVK1L1KY/KIyDqyvT/X7+q0CqdMJKHEhGELZuXYC
EahPcbPPfj2cBXpkTdmGjQE5a2AVGc1Ngf5mZ46sGAGqNQd9jwiK9Be+Am0zTA1e
Gknf83fdewpnf1oUyx5hrHNyFdcheXTQUjbgzNeg72qHfxXn1be8mxpYIpKa5XzT
0xkTXMvG9P2FtuB+r8kj9YXvwy0w5Bc0Hx2ZV00DEGmP2znYglZdj1qkTdyKgUR1
BYPFpcVNwAZB7FmfeJ5daGnToiovzUu3qphYC856CWPnZMRWQboKkgphfJnxetvT
lk2Z6q1K+mWNcFGfh3DTX639kb7kle7czVgc4ZJoC6OB0sTjvJ6/NuCw4THzbfye
VFOpUmX90/rvQhKKcfJ3wIWybdXRlyEEApQ7Jdie7dPM6NI2uDTsYV+FW3K8K2Om
yY2vW4NpQMl8zuyqMw3QKETLJzr74eGLjIoFi6UKqzCZyGpY/nwrga2b8J8jAU+P
QfVZOKl2rR+xJKI+thMCHsaBeU7GWnJlz3nsjUSTIEQRCKyJcjww8RIi92tvY1CF
79l3/ZYDcZDokxtRcjON28PsfuOHOa3S2lelneUTW2KDZJ8z2hk1bzrIB81nWEAK
iaFms0OLAnW7KLC4LVgxtzBpK2eNgMNh0YE1ePWCGhYqsnAit2rBsnyytTmwUGgW
wXEZAz/YvFhm/fgvnUPbSb5f5ty/cE9xDATjhc+qbrel2gFRTJnQWq8/sJZ41vHv
HGgriSFYW51vKunyPXXlKz77I13iw78oL56jIDkVMtDPR5EM5oUpAUb/GQvVCBib
TEvJyJQGfmQwhaOJu2xmsIpaZAm/n5TMTwk7rtNkh56jweKfZzrZfUtZWMiYEj3Y
GTbfVOnInjg/EcAVhDcaSgwoYO0Ln2ks2Vf8X68/rDl0HcYkWU04mug0iGb4hsWL
mMCk60r2uYPxNsVl15UxW+g2xfwk0CeCEQ3+gyHD+ZqOb0Fc/5yxGuzkNHzU781S
+gOIbpNLN/hGO81U7y86qp0i+lmtYuxDlQgMrAGVMEcFzjIH4fdWHeKXpsTvp+nj
vetv+MTvEu/BnGOjzho6LX0xvmVFVgicf616aWKQwluEvFy95beuJdrQWSu2WBwA
U5jmabbVX1CdmNy5IRVXHIfNL7B2sVxPb8qM8iafSg9goqHEBiXwuhPdG9h/Q5bO
r1M4CGe29P8/gJpZ5ErR/Y1WRRviJEpjTY9ORhc4/ZiS5rnF8Xc0uU8aizrpUFeT
0Tyj3cXvpE/hjs5uLqdhIEirVIUTbi8YrrKwuwnx9aSylLcccHNtK8181P5OENRq
dS2d5z5gq/viHYh9Ye0vj83DiP+I0ZEjOYkR63aiKQ4ubDruupKz6PDqRfkFgPIn
rw9MF1tg129zNqGP9ZwztiG/4oZNRCBEePIQ9k8NA0dC5NG4Nqbuvc2WgnmPimWC
gEui+vEx7MaAqf51BFKsnfIM0wiHD0thQBQnYnA2btbT+3LDsNra8d+wLOrmrVy5
IdjBV/t9Pbk19iASvoebzcSB6IQFdlAo0csAPXy5ulln0lT+M8icQg+1k5OpUl8e
5C5frOkaPrbWd+T3ENcsf0EltYIsqylKZ4IAFfjMRijJsi9EvD+m6ZOJDI0Xc6bx
kLVfo4evOYk1AKFgy2RuDa0IN+yQmPa5kfBO40NQh68VfcGArc0sB5Vx0PYBD6sD
ouKFm02xazQoXBbw4xfFgBcl45XRYH60B6Wa2FnOUYwHWAml4H7mgKwogKuszTE4
/KlBLeKCjspqC8mMDXlPIgd5SdMHi9hLDOZhJtew3ehzI5W9Rq3uzHrc7PQTNT+Q
BWb+pXBtpsO0zd+4eCJHXzwDiVTcQ1cnaLreaANzBP6v0LflZVIQWfkihZ1wpCV3
6DsMpS4B6jp3ETR1+YQTRBKP2a3vJiJ1iqif5q7xHFxPNwLT/Ejfok2tNkpsJQG2
tIG/kGee3ganL1Uu+0ZnU9i6g2ZDho9AHKk3rqyJDGOQ4aj84MOCSmI/GsValeI0
pq52EVsfULX/2eRkE22cNRF3EGXu5wz0uematO1RhfSFPUFSMzyX8OXmeWu/09mN
dpIJJwJtK+21PDPskBlWwQ8oSXspgJZXZG7DdAwhbIq4vIkYMFUlX+nIaQ/LOSfa
V9d6Wcreq8pjk3WlQ3WpHrKzoPVzLHz5QLjnGb5c/NyTe/S1fj96snc+IWiQjX+4
AaEMiWjjxS3vqvAvoA1BORuwWzbMQFk7JpCmAfQhdId/LJAZWmAxVDVHCPLZu+b7
UWEJ1AmvWOzQ3VELEekM7bOtKSktKtufT18J3zbTg7iF5cPyT5H87NWgGW78c3M8
TLNl6G976vknsoQIe9suy4Wjb0+jU+zdzaiVV+jfnGoQdRGb7qcQFMbK9KiCjhCl
T6mXc8ehkDuniVIBmujTcC1EM+w/NSgg3Q44vrz5Ku/tEkMshX+zYMASOCm2pAk2
9hTwY8t16Zops0T86KOdMNwHxTAJnypM8jm3P304sQKDx3AtIEoQIYHc3a47EixL
7uD6ZT9M/GO9dRkM2dhstN05js5WSYhffFbc+Ne1RiWlVgg3SalaGY2IkF9Jt1Zu
HIadyweYnnLfeQNBbmTrlsWw8LuWltYF90V0RxQk2M4iu+c/TOctSe408LvFm72s
ARdKIFddcPrNVB73+uq/r+6fevJS3xEigjAn+skwXiNsZCQUhr3e7llXFIcyDOU/
hr1HunD7I4362tExqZpc3B0hZo9SenChWoCwCO5pYBcCvtXUX74n25GwilAU9PPT
UKWaOF2jrMmsD8djDauLie1svK9JV/R28+dEsBWW3OAkY7FuUEU4jzh0E3gXn5pr
LvQxeKDcWLKSC67m6T7qsVOd0Nj1C0jl+WC+DHmfHh0TXoFgEn746lkelsfdY4U0
DdPmlU5MyjifVTr0bEYiyhTO/jw9Fa6DesonLRUMRWWb3UkTvU0q7YHAZASG/5zM
OFesULlWX6Gf1byL6mdCTSPQJr0ZaxxyKgG/YGScoZQY0GaiaBQaclqRujOhQ9tC
kNJah77D6s5GgTx9/iNWLm9yJPDF4Klp4DKdmruP3YkJu77MItWBKo73q1s6cwqB
cDRCrYxRB1CT7xjgJmjCyeGTPKjshfFnPptWO15CmZ48wwD8IsT25XNkWAgI8oLD
zNolBFGmQrDWinZny0oYsX1IQjFxkwFunhvicpeF9p2jF3cAN8uxXfyUbHJeThfn
4GTetorHNtEoUawZQZGMRAHX7colvJejkLrM2goUuhxKLnBlIlu5HzEqqWX89GTR
3kDaeXbhc8OflPl7UXEFyIzL0a5oV/PQUV8xhbL8XYTCfOTONxrBw7O5UU5FIOfW
krhRiJEZj0U/Q99JxewdNEhTUTWdAPHPDxRZ0uXvD+F1zgHEvsldwb8tWJ++mVN1
ltQVZ9AzoPdluVQL8kfBlw/ZMa2tby6og14LKvvlJkPmy+oudJk51sK6CBGOCuUt
3tnkespMwR+Zj/qAftOJOgfhglhGtES6pwiFzWF/lP3GmBiTT2m2I79n9KxpE+SY
vPnupFMv1KVFQlF5PAC3Q4DoSKnWvtTFOEffKzJN7/HE8nfQsm3w84OJTC56BglU
3Dxtg6MjX2GUMo4F283DiN9k4v6yYoBz6BM6uBV5KC6UQV4b/zT28nJKlqHDmIKn
IhQgE4A569EysqFMXrslUb3BtyBxtJ7QdVA2aHqHHHgBoBeyjIsP7dCQfdUr+UFZ
dqB0Do+LB1PcRxTZXSa2+MAB3C2+gOoCShhvDDFxpT35l2UKm+A2a1xKJxXog9eX
o7K8k+/MxymvOeyVram5abuuE3AtgOsn0C6bjvnzDfv8Nk0BWm4NahLhXYAOIxLE
Xv9CbUalnZce65qVvWoTx28P1BEI3ofoHo8lLtfoxckBGBGJhG0xWGslsF3qpScG
7inb3ZqzbKLbmJVDiCrFuNBHUgb78Ah9yRurvND0xNJBM06mmZnXqfrZrzMwb1JF
zRrTpJFr7t+r5VoJTeRpijgkRH0YKq57hTCDhH799XomaXFbJ5S0lDtZW9l0OJNO
cEHBf0x9JFof1xE4zWLQ8HaeTTDLM8LCCTFnPbY4LNBeE/yukTSGQ5HDobEX03Nd
C7PUnTLi640Fdsi4qElillkyTApdbkb/L+JXqc0tldRRVgiyUvv+5SjKxOhb1/aO
jDpt6IgGAoM+TSZgF5A3G9zHUZu4wwEJzrb0sCNxLAo1KGmy7FfGFawMRYsBzESk
/hocwknj1z0t3XoSLwEixupp0bNvYzOF6NWAkmKpiY0t3icFof9RHBlsSjP1ShTs
mEk6BGzEux+ZYJ4QUeg4TZJXOnFp54AR+8xmel/dgWIzN6qUjT6CDa/JiCafYlRb
R3aDAnn/q6D0cMMm0Kzg+4+VN46HA4S+59liLazqFhpTSUgviPTzt/6hMjXMFCx5
Lq+igiMakph0kdwewT16jogfHiJTzR5gmtX3kirBtxL3FTSzTX3QxgNJJBpEOoSw
7FJ8EiKummQo6iNI5WTk2sgxrnG/3DcGpR6+fOWb0hH/Iq8Juga8vqLGYQaXSb1V
wX1IeGCM7aPZdO2/BGktI2XTA1FfB1XQHjglFF0xAqRZ1GLo+wmOMg4MBJfq2uEG
6zxWquY+8/joEaV3IXCLEif7OSRwPnkPEPiczX/6vE+ATFHb0VX7ub1dsfZ3oe1u
BR9z1EAKMJ2HbTEg/ZwGFuA5qHstFy9YxFd2h2PdNm/gdCiikgx9iEtzVztKXNSD
0/dPVevEOD86WfsG6dDzKGie8Y6HrE9BUUlYg1UjPl1EwADdG7tskZ8oY1unPNGM
1q66+aiFC/oPOdTkgxLHIcyoa7ExBBETbg1qf1cqmjmvMQJbujfXQzfMJss17DkV
T8CL/5a0aAClaBnfNTVU6ireBF3SRVqVCnRJWWeK4SdSCfcay0w3nG3umxhCm0M2
EumZF3RQ064uyU/9k9+c7vEn/rMcnroEjVgW0QIV2L3RWcxFeBTqzPxuQrm6vNyc
vAjJ/SffYtPKfZ/Z6Xcsqh7pY8SjqN0Qx65A8O0Iq/abop90ouTHxR+CkpIgsmKn
9f0my1Ti62TXsFuAEdOqTmm/XFggYJ3V6AIFqO1ppXH7+OP/RfgJF4eARh/aZML3
+WKPWJlC1jW08vhY0R9gxVGZNqtviUlmTOgxI7dh5dRFvglH0iY+NX7jLQAnuBY0
npzAq9YR+yIRNiiHj6oqE1aN8VZqPNOXlpI2VbpV9Up2JuJTbqzTcCZ7SY9SVnTK
l5jmtOZo8OnPq/GIWHW5eS+JB+fMmK7tLtvduKgpmADYOZU8/sLNAtMlqwkMNDMA
jEZKSmFFQrVg3dLk0Yi78koihuLWkPynOYhX5a3zj+whIdCn785DZ3jBh66Ytq6N
/VHXQkA9yiTuf+lqn5ZHV+ToeDk+khBgty4kbkbW74qg1S73HJlIHR4V7AG+dJve
o+FRU/QINF2DU82ZC38MGNyN6u5mthOWq/Ffy5zzqjLNOVNQvTh7A3thmlEP/+jd
OjoeoxQ8pxh4B+Qm2RG4NXDHgKJcOOHvjoErWicPRugaeMthci67BOq2S0OxjIUQ
QNiIMuoLxATQXtTbpQskuSFYfttfQCnGfEI9ha3Ud+H5k+UEY3nmA7W/NmmPMHCR
370QVDgqAT6SrwtFXONmGxCu9RKYPiLALQm5WG8fUf5pVyP/HhGRSLkHrb6I5wlt
fFKj23irWzuEP2t3jOqKBMc+9eHjMwXJwlEXE/dYEI7+C4rxsD6/3MFZa1QSD3Rj
iweiXM/G7dUjM2fPR0RSfMHQofmIRcjiRf9nCQ2HLFeh24GtG8DPUwItP5ObfDmz
xe9zuVPv/NNxidZNyxDM3VZYqSiR/L9/EElVQd56GTOgS3ObyHfJ7pyBZxPHJLTr
rmJS0xpN/YF52xfz6IjqwoHthDdsjUpahdMrt4hVYgYCR+vWsU8szADBgPxjpVQl
VapUNxC8AmvPZVXkkeFM1iXarht33lf/l7Y0jgHtoi/B7oKbn7Gqsc5d9izviKlX
J4uhTXxrv1p/eys3q/mCC4y/YChdaX2/ziEpWAk0BD/FJk2ln1HlAdTUrBUeKG4D
kaX1JRG/3mQv8Ps76+8Wi6mQtS2OSGslPHBooG1RCX9m4UBpQmYkh/68C7aVkH7m
I7ASWW2x1Z3Pd/IHAJturfaO/WsJheCoYDGhJnGIucjZWHdcAwF3zrPeq7nTjJUb
UhMQETUzDPjLeIVw4j1itF2NFL5iM65DvuISTHZPuKFzh9DolmsyuWjO03cqnsZa
e3T66EBSu2uOxpb2w0IenqcpbQLVz1OFdQady6M5WRjKcp1l7KS5KdWVn7NmTkUi
6/pO8ksDfAvATLBWentckpJrSvg+Lg+A075qpx/PKDIfP+Aq4MpB5nmfULR90qnd
RQmlgHtRIVKwUJQCTo2C6le3KWycxF6j9Uo9nIpgwUPuNWXlKdpe45ubSDQwp9+i
IitWL05ok4uGlCRI0elj/lxiPc3IhTTa93VRaSpt8TOeEwXXKWC+G+7iriYbRWzQ
S2junqYHf3afqoIxEfb2tNoq1XrTgwLf3oSdREG5GE11B6dDBiH6y6XrXTCJ+b3D
buPGej9A7eo6uDcPz3X0XRhaanhKAoFHf46gRv3OB9/LChUoQudzV4Q9655UrPZZ
b8tkJ0R7aaFBTVq1G8XYZThz3UKdurqfTiCUlWEXL+rpS55Xf2/os95HhMFa3GcM
npdaen3XacCPDtaaQkKLsLRw1d2niVs0Tfm+gTCqMYQlCbG5QjIp/EleXte0FQ3F
DO1C3k5lcGHe1ZsLH3B5XzyoPIDQnEA2nfVEVcqcw4PBE9oPl9n+TRwXSazulAmt
gcrFtf464HRr8af4niuv3GGOdL7A3aj5ccJ0nB5tybU6k8d9vG62p4Szv+OQANzQ
R5WTr3gUH+ADkPhor2cNkQQbtXTtCykqvTknA4T/nuVy+Y2Rv30x69AWNCnssEos
QWizQQBrJoKLPOyLkaozM3fxRQM98Y8ekMaWP3s1VlxCX1X6KuhpohrgznqGTitA
TgE6KiDLNRtfxUYLYIMIsRu5W6VNWsbgPzaz/OGJunjkQQC0g3APME0R0/pgLEGO
NbLAe6rbX/vkNxNEZN6vSvWXav1J/PybvfuVrBeGcfq58FNjY5hx7v5LDtxnNmnp
8+8F8TzpYq+l4f/EeT1nhCpmWa4r2ORt8bI5xaXlBASUCy0E2SYoJXcz+PHKIc4f
piBUMmm20ELtJE1r+kijSa5c08tw5v6LjINLwJcrbcBx1bu9Kytz5TvTWZA29ORb
vQFVF0yOLWXYDzZ5TvGsDxfz04Pgi4x6FcFkkOvCordRGtKm6PkDnHrgwymIibYl
bwnWibQhytYE1v/upBE19KyO0sml3ZXL9jMRTxzgzuuKUEcD4RXZ20eO1y3JnVDf
oxUTvj/grtcpKp6NvJAovIU/nrh/EvTH3rMePnFaPv6in4O8I39oHbWfawxrEwCG
aZtWD3FLE+51FO6k9VNtVCLS7FzQV3T2yZlzD0D6G2pI1s2+12rO2eEc+s7BRuhJ
GZi4eEeP1FziE88SvB/WREwaz0Rl91pO7HP/djzTrWZjKSf6rDAFhkWXd3w9MShe
xjSUzo3qc/ExvDnYbPxoBKFkMXt1QbePFsa5hU/YybV8VvE8VUmatSUaCvYhekaW
XI51UiiL8F0lemk9O9Yv63DjKdGOvrT1MD2Anj8sysR/1TvFGBOaHG/dY1WXhcS+
OOoCrMh4ZuRT9Ezl9/yERoUuOvqw8e82uul67Cnpm8rm1BBCiANXCnFqFq+0IBHe
8Pnry02owAsQEq8oP3Nh7T9rm8jarF6dB6h11DVXe0w47ip+tJqW4LP1ybXmJNVe
e1xe6iZxMnFgsesvAsHvx3YvvEb8P6aDQUg8yYJbji+jA36ASflFOREFZV8SJkRd
La4y5NN1ldEjND+EF+CavzAumqm8axEqk4UW8ThEFt6GD2TCMBEN4EFaamZmjQaf
mrTRBzAQcW6whN6fB0XMJvVsYq35XdD+CIFTxLxztLIPVr0gVxQVFzwBNQi1v9rZ
hMA1cJFVaQj+6Tko/D5aYyH8PkOCfN56yM9yJO5i9s4uYtJPZupSO8O16WpDFX7Z
pVZb3/QboZcOHsXsyDbhN7cjBlhx5x+/5R2VnZYyEp6J10pYT55Yo0zD81kxuo9K
zSQfl/uquYj9baMYcYYrW6CJURX54LSuoX5hADs1K1obOQoP3xraDlvZ+pT6hGMR
CuQM/xerWX2aqwvtk0JuBoFdEIi8R5oulbqyT5Xrkr3mr17YfoHp5zaz2LUE+858
H3vYw26NVxZawAdfEQFo8sQs+dEtIYStjIs5CF43YuzbvoxfHxFpidOaANgkz+3J
5t/zizl/VWOKY/C0qB88SgygcJlaIxsMBGh34QL5LDo=
`protect END_PROTECTED
