`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6H3WdRubdeeQQS/DqJgRwGAyiJ39xw52ynKthrAENUIdX2k2aqy2ZvcINSBMhAyU
cYyki3F8ubV6HV+a4lqLz/XQlLoXOhGwB7sKFQpKxhblk9Mx6sVXbKY5Bpn8d9W1
gvd2YuZAtnKGZyx/gWWRAlmugbrakg6KK3kT56FSlNgOGkZB7GQUoKqxC+k//5hJ
/B7uEugLRNygW/cCHt8pClJW4P5+6sXR5IZIri5KH3r/San1VP1NpkirSUEf49mZ
1T8SwsEvOkBF5WXirZmulsoWDMcLgrN+ESiX5L6IJrMo4zTWRKPLuxEMH/kzg7Hm
fCkp16bcVmK0FO4c3uxoVodIgIcoOR2ND22JY3Et+XH9XZgoNmqV139t6/amLxnl
OweUl3j1wika4vNGfAy5l9cqPlfj5Z8kXlyUTNM7ZsTd5es53jjZS/xHTOBUDf4m
BboHoCyA7RFZdGlpyHojxtyDYhb61MGsNfSe9gCfYTJKhzHmS7mqnnO8hIknD32/
Ak9J1oLVFWoyEH7xQwxCCaMswQ/cXhDrJ7sxgCoQSmMIacD1D/YG2g4dK/1aYmws
GhUjKP3A9xuwrqfVxqlvC7WpedL3gdo3V1M8hY3edmhVo+YPI3vLjAvxcHrvqaCp
CBR4hFSqXrwEv6/NhvBYEA/Md2PIJZcZByU6ZOIIMj34eNWQe5JVb1kg+WGeWMlQ
B4vFXJY5Av7C7S7er19tC7+nwgeWX9l6DV9DMltjWav6oZ1irzQuw9pLW9m3zstH
Gnhcvvl4dzPBcsgt/tgYnsNjwi2SABY64h10zx2+GY2lkjYg2CusXIzbInmrslFF
zkr9WTQVRB8i8Ck2mSSgetjzIjvACVLhLHCKXKhEJh+s81zZIpTJYIVv6eYp/ash
ayI8ULNwQnBM6k956/bVh7G1OvQt+DirXN/3XoBngoQG/SCO8bXCAgO9ajR1UagL
6scsjd9v0bcsQDeCca7lVDm4LlxbRMa3tMQsr6/ihkitM0UYhh+C+6miA7U6/QMo
OR23ihSVFR/mME8AAUuQQ6P77OZj40jaPxWDdZ/PTU119iTywuuMOWF4LKVqfXpD
6HMjcNVmRAEkDMqM2u17l69EmgEFUw56hkkL/yKX9ZLMAAco4pVv7GEJvtvi9hjB
y9X9X2jcS7UU4HEtUaQB6hLHZhMMzBZELaIUPQM7Fte1OaGwN/H08s9xjrWEw4Z+
1D5Who004lzB3us+yM5/1JNuljLyvaf4xVatYYjXibKH1CD1WFQ3UEH2X7LoNdQf
DZWsJ6iimveZQD5nZDxtQPx3D8VQnXwClXb56xzxZgssdB4Fn+0NxXRGbZymce+Y
eRKzNM+5znQ4AsQm4Wh0VwkJrBeOtDPtjAWp1TK//8RebVVsYp6WnII9euH8Fpgt
s4PGsOLWDj2oUoa9xtEIuAzopZhSK/V37PD0mO9agy4ELE3aFbC5mM7FzHYoVmSs
WxzhoFEg5nuX+y4b2yhdAiHRMhYF8+Z+UksuFDMGTIdwxAhd6UgWLq3ZkG8GYIKU
XFq4EvOVDnCuxnejM6nd2qsFtjDE8pjUy27koXBPhU+1NI8Zs0/gBmXwY/rucVQD
ZLVdRqAA3ykhZgKslcxDnhwmpOFgxia3QkeGPPRtnbsh20ZinACPYDERzBY1Zj/e
hNHido///t5DZx1z5fBcX7Eh3jY2+BEMDLN5nJEI2bOBdFkai0w/mrexDb1oZMVT
hLid4K7xFzsVgaZ7I3X8KVuDe8I81ISW9HY6TtDFBF1z7O8rxtzANlio/s2soSLq
OPiewvJ/NoW35vyneKCZGdUSiuP/JpY4xrO4o1M3MM6sEezaGqCpODARHyINPqYS
8yBcKyMqp0DTSrpXTfwIzwE7X8whziuuukB0PvHaQ5Hyya708V4TzWINTztuHum/
SeSjiyqUmi/WomOpXM0kLSHKdHo9/7bzEJFNesRp4R4+JnnTbqKGIVyROGFjeIRZ
GBuTpuLEnTFse5ZDlGEe7xWQPTAuQr6JRUp6xTeTukoPydxxfMevd0halxHUPtbm
6NkPXj9W7GEsKiTBXaZL6NTcOHq1XftK3uJe/5KYJbFuKSrlNF/bwQDJScr5ahlJ
DHYi4GnmcopYwImSzFZRY976rcSUA6Q4GoqIz17b2W5yOwGHxQy7lQdBCZrXA8At
1S+IjHON72oe61c3j+DdC7hKgLUXAze9Rix2MAuFp8TRFTaBhmb+bUHSklmB7Trn
+/HJ9E7cnLaSsrsqGoMSM91kkQoJAwUVoFDbtvN5aSjJy+8PofNUJ5jEvWdenrg+
dzjTIySvc8PbLURJUTvviuFWbsEG6pkiVGi95jZ/Y9Es4lU9ONI9xf9DELY5UeOL
qTV4ABW33+vQUZqOKeUx4ffiRc8MRZD6GwISa8Xf/iJGS5ymoW6/oSSxlpSkvZLu
TwWNeEj5bzZfXF+GwnlcfhqwfW5nub3bIw1WSj3pDzSP+r1G/oD3cWuW//ASNY02
nh4d9I3qGloFNbWoaxCXKfq3xT6Tyuky1WeIoMAaVomtJTCKwFABnkr0kf2ZV2UY
yN09MzLIUZauipDJ/sMkiRPPuolmWKnL0ypLza1nxkpF/8MvnPQ7GVnv/c1O/P0j
mbSdYqvTj1x2r/gzpmI+pnXF5rk7MRdc2pCQhuSZuqXqtI7PSVdREmQsazF3Ix1z
ZvVkX5tFrNPK6NB7MKCuQswydKqCdS9BDs/7X69h18gBZ+KRBMLiJPmROD4CN0ot
yvQFdo+slpB4VmbEMKTlsixOdDJ7whYkSei9fDyMyC56gamMAo9KQLPtpukoBpG6
2T50JhskoQbapLkQj8fU3oNTC7zCR/Mf0mfAYtyC3NWSVEosdFlthopx7U9DDuNK
69Lr4TNq+v3LrRn7Oz/ZP73qDak0XK+kCYuxlO0siEZj2eqX0db/p+zVpKxzVsMu
JGNrbTj6Gp67AwNjOW0MnYx8LIorTLiMR68amqoWgV9cRZTUL8OfSu1KiZYmUgBE
owWXF49Z/KYxo/XUSs64F7g8EZNDO3fAExSrcfcry8fFgCZ6ko2iqlqzb3uJfUoI
3T7sGhVFNAN6oxuyLBX+bE7Wozn3gWCrSQwIYEvqADoavhY6PRQyME4dkm+VwQE/
v41pGgQY44qD9iiJnKjBrv+pEaZBlvxuJlyAcPu4dDSp/kMVOor6PxxPK2iTZdeQ
UTi/W/YI85M1mj0Q6ipAFgVFKmSMh1bU8jdJvbMUaMD+CETfIjBUdm+76kU5O/Ql
n7axGuCGDPusxZHYkm5+T2rSFqm6Uak4kgNkALtJ28DElqecVW4ZndttBcCkbJlG
mKHDWVq/Mc/WvLmQZJCg2GflcrWBZ+E/LLnnbH3FvbSOyf0Rg4sEcMsLpOi1dgSM
r5mYeeYCvs6RdzHYA1eZp6bHvU4nXvHV+4EhHQSAmx820fAaB7GP/fQfQmXiyxH8
e73KYDsx1iZz5umGQ4gt6Hcwl5Orj45yc5Wmkc9ykE0ozfh9OJ+MFZ9IHl7h5c+Q
+1LHHxSa8R3EZPn+oNvQ2JAkhsn1Ozo/f+mIY8yUVuTFqm94efVcwPi8+p+by9/N
3v1wlhVsJwtT5Ys0uoBHomoZ3LoCgcgvDt/LvlSybmt7pxOzM5MkYdCEr6yefR/M
S/yR2Ycv0yn+q8ogYMQGV+b+6w/HHRQ9q2Iw2u36yd42uS8leqZhHkHXP1v9oBtA
2ZEJurShkt+fr1Waq3FHOlYDfsxChGS5SrMPZXTE11+AORouca33McGo8oQSbZl3
VfPDmxr54N7X2euMQA6TOAfDhGNxSUVqdBaScTzrFteOABmtBGj9WE+e/1ROulag
fZeP0O6KxwOZZGX1braBkwrJqLnrVsAawbQ3fl4CF3b/CrxFHiKu5qmM6vCmwq6u
tqvjXHT64Qac4AC1YCdUkCbV3VVK8Oiix1yNR7/BR3XjqLTbzBtJvOt/FNm5UVDL
y2Ix8Ckd69aweS3SZssGwSCqukog98isBr+naDP09OW65HiYX9FtkBRVezzKC7zE
N48h+Iwbd1zicjOEhuo6dJnp0ylJoMEVcbPZRNTGTZnBj9eDNH8Gr5OkGfrnC98H
G7Ayng9LV/93EZXrWF4cFz9WCOYJMLDQTaiHT19GcvANJMtHmpKZQZHqMuo6Uyk4
hXZDdfHjqcQALvvDmVRqwzyiqFe04/bG00ByxxCXSqeG/HahYiRXe1O7/35ODQmZ
/3nLm0GLJr/mlLRVZM/TgdVeP46YikNphqmALjiVUL+xwAag/44Txg9GALy9L/qk
2b7tOWSIj0IT2cXWS5uDUq9lTR0Qzg3VlQ8nNDF+KH90evWzwpaIQ/4C4rdV8bTf
mSMQGOPgAJD+06eCR0ftEVt+2OhM8xql7jtd+Xobu27JSJ0lxqP4RJ514zW31tM1
reM6CQiHeM7dst5RS/pac1QYsaWeBxQ89O9tricudJWRet5ljN00rgWyDHGKXBwj
gjwb2JJYP4HMFq5oVGPn3uZwxowdwQBdLiYMNA4YVlD3p5dMWG3Ct92f9IYLEZt1
AUU75TO85AZNPY8tCWFAXc4C0rzHnLQWWQSBCZvfxCmY49CDQ8CfpzoAKTKL/Xk6
zFfPVAUPH5yglxQfi7DKUcD4DFpHT1+nG7RYf0w6YMOP2Pzgqv5OMZXFDQMmUOU3
rA+tZ3g5cReebwa/biZgpxhntnyKsqNf+muZINLWmrEqPZ4v2PrPKOyfxXNd97tN
/06qRTKCt+qO8hSznBtfZyNcz1iUrXOrHhD/TjcYCOBCEg1LtB0WWBXbnETcAyal
6cTdBkQ20X6gfdoUc7IGTzoBbLltYQvSlsLLHLaF2Dbdb/LgZxgGcI5+YbIzIv55
hEx8CKtz0oduyjbMzGlJOx/wzA19HRdbq/t7yGNsEfPUjiPLXZiY1i36i0Ot3R7V
UxLeEeXaDK6XA99nH4FPwhNYVBy3OQl9bzoJtniWvA/VlJDNdKNQ98XqaRYS3+kQ
ZhaDV3Md0SVzPaSxdagNIlCx4GgJL/KTJUUjCAvNnnlj6PeI03j5wjl2G+dwfTJa
FvrTzIGswfmrNBH8Gkrlt8NPuCxPS8pKTmrb1eLCh00+tgE53B7FqxtFw8FEW5tJ
stz2ur1zS5lXcX4NGZqCPLKmcGLGvgan/DTBwdQua9szqb3zOV2L3Q2wWCoR/5En
E2VYWt/nLA9ItKgL21sviXUKIuvJ+KjR3j/8zm50pkFr0wWZQyl7SnsSGbfRpDZG
rOZmiLGrmAfx62sX37IcAr5Iipp4Gja32EMi9nns1NmPZ7DEeiymKJyTFYZmOwI+
wcYFHCURB4lpirtWbRcU7vND6OPcLeu5T95GubnJpbwA39lRmz937axW61Cs0u+S
UrXzjy5v4A5a5aSpYriBeJpB2hneqPMYda8QbCuaaT4NEiId3QMURPgM8OkvQi7E
+NtGWmD+Vpp7PGcT9WJv/HGLrxPvJNlFyXLSgSMTVOsrsinUt7XgzUBulLhduOaP
zximXY46wI5wxO2OzCZ7iu5L+R/t1sQRaIoIcMwVxWAxlXLd+HN4sxFmuOZUdjzc
4uqLh0kudxdUrUW12yBbnRmQioC3rCGRA7UWkdfT/Nak5iOXbrC9YQ5rxBiV4BA2
Ot3PvS4wbxKJOCLpfRaYQ7JpWLcOHzKizPsAn1yEUORL1mq4W58gyStMq27bI2lw
OHMii5K3JT+Fk+0wUYM239aRaN/rHEsORAV+fDInhj2cijIJvazM/8rfDAPFouTl
nYhl5qlT/6Gvj19XMePBXhjKOEqKVJwbRAeY6QY4UQtxxt9H4wJUSo1F/lFrfPLP
gcmJaJ5qgNzQnOBwZeVumCOZ5MlnjBL4rVdyXx5xWD8zIZvcKKCjdzqLKCCwwZPV
qOrdQ/nBeWdmbeAQd57O7b9JBXsQOPbfC+Ig8MqtXIQ8MCKRmipmhP5BJQe5x3Hj
I322YdR3du/2HTKJDgQdGVh1wrN3Uea5Mckb92yCymFZhw+VXwXZIH+eFBUycrxN
IF9usfvzj5ESYcvzgmXTol38GK0V8GwKKLTEK7L6kn33vsotMFWkFBvefHQU5Q+5
KRBrN2u7ZUPMEuo2cdNHwWzGxO3sNK/+2y8vBmu0ksAb+BkT4cpzs3iSXHJTi0KX
zB8/AePV249+y1gATMn+6phpubsJrknDceghNV5B4uxzvUqt9ODgNE6KO0tNVEZN
eBuBV/oW9TnRtFxnzrbl3yWas9SfnxJayIL5yFwOHXzfKjZTscsN9nnvB76OTTlv
dHaRuexTJifOMN0l/DPRc6pK1K3VK0FdoapiejLcxD6mr77k58mlB/zcbMyAqz7Y
p4wkK4aWqrxVdTEOyY9CGjmiRNDXwL1ZL4V2hKcLT+ksiZaUuGi8qAhDcSvtnO84
lqUGr9YVhZg2iC5aZMHoWq8umMm1XUepHqVq8IzDtz7NV1VqaS6OlhiRofddsdfY
u34vqDz86VLt4zio1sluKsMb9+u9eM9/dEwubuVixWz6G+czkqRfXiGeK2upQkXH
HfWLxn23dnTyHRMqn27rKrERsSA5d+SZD8cHXut57DzDzO7+RGrh7pOgiR9klDPF
qLP39JX8JU/LMCdIh0OuAsCaLVhazyaTURS2PmzucvHLB5Zt/vu8DlVpDZyW0dJx
M1gHnBSr0YwoirYUcZ86yU0YGw7R7Qs+YXddg0HU70NaQAoshAdt5bGwR63Frug4
OS143siLb5mQU9rZQaawLeT5503rnR9mCByB7i0KR+1wYIZR6oGDd//d9q1+qjen
2xaD0FWbuhcUfu/jyYXyd5WS4pW8/0/ZS3Vm/qsjFPYyedlqV6Z8P9QtQTbnKpOz
UrnF8lFtWScff1+G8/Ea4ZomVMZXggnRTPYvLvRgAFRqdugoEZDZl+xMUNnUFsiH
4M+wetFy5iACjzwwexWoHfz8Pvu+XtQj5/8t0e2XLbgWZaeUUv7wx6BSSiCTmsh9
geqRNWI0dMrd5YRTYuDZhtYjEexhyLu7n3cHZXZ+DXTD00Mk/nAsxRYJKWyaRr2s
Q6tOP39ZX0R1rfJSr9hiW1yr1eNaDymlZu+/RMm2SOenFl16UzS1euUMUmE8BKp6
w1rIgorjFT7tMrpkIsntbxvru21lnuoZVO0GmZGPXeV7dvFlau7zr4y7E9LTAXdi
plcxOGnmQgGU6vCO1AOEfYYn5mjZSxWAXqG3bhuVPem8W5XZcyh7mtk6TJPnvqNf
u8vlGi2DWnbSbEHJjktYrLR4K/rnNSK2HiNFC1rygBA0Do7yF5qfOffJdzwNWMnz
nDIcXhXAOWWdpC6gPYhG53dsM43LgYPZSqw2dJYnEGe1SR1MfT2s/lB1psiDvmUC
UmB1xYSWItnWppc544SIofTFxNrw8fWZqnkdijg/WRFFesPgg8jr/xUiui+WWsbp
KReQRlSISEPE9UqtO6fMuvju8d7yNWnhnQppM0/HkKovIncgfKuk4wwLDS/gg9Bq
EJzdhTFXIrR6TZhcA/uPL5+7MwmO+jQZI3CxFU+YC1q5LOdxwNzweR1CdO/2eez2
osbnVA6c1SFKbdge/HQvGq98Ii7BQ6148+nfldD8SVCN4kZROZWY8LesOkqkm4K3
s3isjLAnw7GOnVDlY26NeXd4OQUw1sqK3g4xEPE//mMxml921A7wne+c4PECIfro
mMuLPoP8izfDS6CGkgpI4PSKzpBBAQCka1eJ6YWrhCKOLYPGo5OXq5kOfXDx1gFC
Z1kP4rwm0mT3tYNbii5ukq2fFoc2+31DlSahsXylEnRjVHE3rED5Q1a5RRxsDyrp
u/33+HEuhX3GtQpx0EpZr4WBuIRyYFA0CN+iddrzXUKjq3KuSlZhJM1Z5UV8iqih
dYXxyHIY/VwbgJe1d1C8oOmrPOwa0tThicBgCkExI5bUYHj8cdGf2ddk0S+HqMKx
NOC2z7Et9lfndzJcYWdG+UU+Sx5af8tcZLxCbNdmhHeajSoTuOweQFcuFpgDasFV
nvU/vxqMZY1RTEjswR/OaVS5/vprrkNH7I48HASfW0ELYYTZcpC25EnCCyTF8MOz
MpmjS9VkDdkymvsjgSq6M+kr4Qi2IOtNzSFX2zZ+YSHQv1msPZptBKenwOo4gbKj
IXdUb3ZaZKeNznKMfaY6D5pAtyR2HFa5gabI59tWN+CWFRjpMxV7GEBgNQadCTL+
UXlEIYR5U8voDg/hNO4vA5rmOMkHkhzHnLcdFXxNKJNriVZaPxmHW+wEc2JSsufS
ZBy2V+4m0PWRUw1AE133pw7rBq7nqtDlKBKFRgQCTK8T6uBrl2UsY+mnIRBG1RMY
/Z2SKCw6TAgdKfP8o5ugMMpxJKbKnD3xmAo5hbKVTehmIlsx6kn8bb0m7/AhVQgZ
W6Zv31t61aTnLCu1ekNsSRfbLfv7nG/pPSWf4DD84qu0uasW2gAx7xqDGatOVyGg
zsSJqR1I5fSv4fIhut56dQ9NftHFqTLxFhxh2iSlATMomQId4n2SaSjSI2G8gQI6
1mVHMkaFf08cnE0Y/aYX3HH4ZMiLK8/QunMzDQtJaCKIClJFMr+NNQ43Utnn59ZS
0ahT9UDaRmGNAhwQ/jhQjfjlXkPMz4GszZX3chc6Fyex9jXjn3voxsCB+Ilfg0cQ
Vur5qwTO4o7gyIQlHVJY5j8GnS4gZajLUGHmUtPx2zSeS/1JHP8zQ62xN9wItKOK
Unq94KqCBZuUxrQW4F3LGwCSk9wzcEJBfCsFaDU+owZ882IZkVN7GwBbNwVaFG3o
UoCNcSDdCFCrGV/JxbARlH6ylParEod5wsu7PN6VKLAI6v5WYi2qLT2XRHy8/G4U
9505QFJXSIPY2zjNhCUh0iPpqTwMoAVziCnHE6SrCLQCkrYRwe+yExB9fZlm7niJ
Cj3+4YPd/i28mpC4Q+H+knKS9cQF815qRF5ESp4MW7k=
`protect END_PROTECTED
