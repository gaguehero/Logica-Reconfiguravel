`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hy3h/y7hvJ5jOZL/Hpt2XhmUPS3E3BpgalcZP3x+B2zF4ToWmU6Djj+Jr82ah+ic
Ei98P5UuUgdlOGmcqaJhhOROvetLEh//RwjNNCR7IdqDuFX0GCHOeaK45h9cemEP
qE77mYCcls3ta3Hj4TK0m8pExR/mSNyYI9+3NajYn00bPCAoARUlpl2MckMJZ//o
yIp3n4qR+R+zEt1u8jfoiGXTlVmDhXZ+LBj9On2WeahKigIXk8wV2rhW7eBIhkx9
+cVd1rkJ/Z8Vs9t84QvlAEyTOelo9w4zlUU40TYno3Su6Zdt47lx13GZ5IItIMeE
+9dlGXXKP8xBBF7p5G0lyI2qkMe4/uwTZURlIdG0fLMw/jVtHXO7HhWWxjOMaVR8
EiuQ2G23lgxWpODNzk9mk1DDbkc6VCHxU7uYYflrsUnqSxdjt2jU7Cy+JgOxGygf
5mhXo1GKt34WyvI4yyEmpZci0xdMvx/t2KuFqZPG5hN6KirHCr5Q+86IhRu61Nzu
g5YPxRn/V30UPp76goT2AjtXJuPH35o7hvnCND7e2CMNTm/5NgOeyt8P2z0+4B+u
uJwx1sYTuaR2lIxMn6KAKECbpgCt6X6KPikpYMPiqSw0B/uN/5umnClmXbdz6JWf
Q7gEenQD9uSWgX4QJQ9H63egndBSgUMIiHiQEq5swJQZ78oL0X3fDp+DGjjtR69r
iiPUjdrvU3KaB3Z5BZDEaswqgtc5MltUcl5zl5AOaslqK7dDawGf3RJSgcz368gE
0GRIBrMAf0K+TryxLFCWX6q3rkxA8Rvpe3EMyi04DhP3S4mwymOuS5N/hPESj4B/
OMYm3BMiVpsi7XDRTA4kNTek0SeUQaCXcMTpLh5HAFN7YWbGAqJWsJpSWXr3XNOK
Agq7vNuzASGZuzo8eALH8WdagIho/HSAYB1O8Bq75sSF0rU/Cy1MQvACjweAPpfS
bYfFPemTZJ20c2wXgufk6S47GWUMyRl7Fuqi7G3GL1Jvop1fh0H/TKFK/H0Mck+D
A8S8Rg7LEndAResZTUf6JBvGez94dsLv9KmOEtWriyRxbzZOpUF7nNCaSJOXj+V4
kn9W57gN15gjZn4L39g8oeq+qDxeGB+zbZSlRxvqb/FdBItMxEjETkdGGl5W2nHO
ZiTRO1kc7ZC5Qt7LY5Mgc3so8l9Pe816eAOdlEukPX7C8Jln1u4DpDT83dCWWUN3
PV+y2wVV5WeYT4LsI9Se3S+f1SyEY9LOh8XBw/QslknVRp3bpJ2noJcpmP1RTvuM
268JKDxmqEFJk4OkKPo/jkPG35WZnL4ul3F6SyhJ+QW1Zj9J14T9oFwx9bFnSxjf
ucXIMyix+ZjwmN9hPbpnaUcuaJq1S2EqaCw76aafqVmk/765s/YmJxMmLUkcK88p
dxDUWtMA1egEqNkONv8AmOLjBq40MkpSw45uYC+YH61D77PXlZjyTGOXlfoi+9bN
yIEjUJ9DSCQbJ/wxTyAsd06oelvQg+KE32nRWXXek8gHf+iwP1DnXnpY6sSVACI9
Jn6cZydIXoaCwRCBnzkKTA0O+w1MZB/1BaHP6Thb4OsbiUgahtfo2BY9lw9sw/kJ
BD7eCvMnggpfuJZ8HgE6A83HTdU3/K266sWEqJXV9KuBJwpKqtSVMxvk4xjXc6Nv
BwdsD8dcOgvqeqm+yaOz9nfn1uZWVg3zvc9vdtgcTZecpH7GPe6+GE6LlZkhNPIH
bd2lz4gHDYMzAsACa3znYrgNAFNBNWPvM8LMyuqlIcXKnq76/YTRM45xYanqI17Y
Ibi5h5edBLLjdGJb0wKTO2ciTsbIjoJsrU3f1/PdyfO4npX9ahkqQrkoCnLejrpV
X1EuW6CsIKX5P+SL8edlm0Q5jNLXM5fj9lI4XEKngHZ6gjPEd5pUtT26KmXFiCNd
mRZ9s2EBIPYlUbbG1paJPRjn94aanhfS2aK5nUTaJ19FbDhPpAawkl4Ye3wUfC+3
1SAkL3KsXy2nmyg3S7iy+sGH5+QhQx76riAL3SAe+TLw4NLAxZoXE2rziPkNBMuU
3wE83VUWz53/8XmDluS/5w==
`protect END_PROTECTED
