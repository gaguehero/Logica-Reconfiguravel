`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wooozH7t3mxgfFutV7oB43XlLapHxdxNMLPwqY+p/sVmoKXsPQntz0iXGDT0aGP7
LjFoNP9OkHyibPn2L59sVn7QT60E/MC2gMjHtAJsu4BzMrQceUQNtV52RlT3agjM
bBb8c6btdoH6MS+gFqLNn+DCWAITrbCiC3Z3XviQPzEPjjyQAxUuG2KU4tNjFqfE
kUuuGceMD7rkI+ZuaY/oTlW1bctFE9VCHffsohJ7V/jGTIPIIV86svdGl+poQ9qR
F/jYRV1c+n3DMyB+w7kkbYN/D0kdrGyMg9Yz8Wl5qGaVvFYAie/60RjzJDu8+eev
XCXsaT6kL092vjFERh+8XaQoVpIbCr+3CsZnfUko7oHLL8CRgLoljy1dR7QETHDJ
/t9GFsok9yO/sg39MlzG/r8eyTwLZrl8oCkVv/HCmhfDSjXBPIi5sjzTkJZixQV1
zjoXr5hj8fenYD6hibJEC4dqTUPifG/JUF+YkF0W3qsGm/D5j0uYRUq+XyfkARox
J5Z7EO9mBDm0U2ef3z6Yx3dQqLf8lf5sypnp/NrLdyguOU4ojgk86K6QwG6XIqEV
Q7GGhB9yq52gKZDGoFOeQ5Ls5JfPf3dX04VwQulyj2Eys4FUp7rQj8lBU6Ttv4bR
VasyGIcYeOQsuvVR4MeXv2z2PkCidy6KCgCNFI7zxNUZu26hKxb5suEsMX6EMojf
WBgFd80joBGHIpLGCMB2rWl5XLbUKMdzT4r4xDpKbdt3e2nxL5oX9JEe1pN4CU91
afiK0z8Apoh98XvXc1zHH7jmZJE3pEN1XreYdu/CaAP4HYaG6/sX6xchVTSi6VdD
W2mh+aMl5uEqfGuaaGUhYs0zUkbYp/DPVt2eSHAG7exV5w8XQTQAZmvJ37+J39cF
xM5N/BzoYMC39dcW8PPKmaMHQgwlPIzClaxbwd5T5+/Q/lfxh9jjotYJyy5Dg8xl
jAbwHqIdYq9KysxwLFyDXbdD/Zc3SS2cazLKG4r+SvP3eqQGrtr6gYVY+29aRhOB
GW1dHTFeBCXl7jlgy7dtjs4pcDpmoDSQWxtIepeLO5avJ8KfLfAk/G38LZserYBK
XfLqHWLodZaQPJ+xTnC4w76+bpGZOWQJtvu6sSNHCOFFtydSVM+bUdEkYeVRCnKg
LusJuweKt2xPFZ8T8Pus55Mqhw+Sf5+HlGo3GVBTQ/UhIxV4rIq4q5xrCEZ3g98o
vaSv6+Ab3cC4755EMRMk0sKEpvdK2f1VzSo7WCjAEWZI8Q4WhKGWRwO38YE3rt6W
pGI35mC4ouEhsklf9m3tecLRMtLbEbBFqiOdQoZuBLU7Cbo0ZSak+W1CEYnqjzTI
TpS9zspnpdonPb3z9Dkd3n9xGPTRr8YfK3YcGa2+HiO+VKj3OGmY2uHQNrYQueD6
cNbGJRDCIiUYVqpDrif9RL0jv3t9a1Q24z1nfu4unujfaae9npx/IZcJUKk1uSmX
YAN8vJB37IISMMWEJgg1h9FNDYUO3BofLqQqbaFcFiBqR6QHemGTiy8yx/DPISha
wqaUjNBc7yYbEEGFLTs2blILuQBhvp1LIqV7R3/Dyai1dSh6g8YDxGonv2OWLw/c
u48oSSJODrDYaPEUBkJ+Tt7I0ZzaER578SdwaATZABp2aKgwCqNq+5rjfnFSYSBQ
4Q2KM7W5XVKslXZ7EnUaI3GPmffqAjbxqaAK0V6EbOPuGzA9SaqGq/CmkZuYleeg
DNi4/9+gHT/4g8PEhZmLzXpkrxJ96fh2Ftp4Bkx6aL8JnOMjr/9iLgt8+CcktUQm
kkZk0RtQZDN2q2CAlKgfBdW57mAuiyxPcO3v55ReGIZuQ0WR98BJlqoX+A6OLQhk
wOsDd2Q362eDE+hs1qZfefH/nk6xHNQg8FZUNXoHR7m+vWlCH/ANVabHMAwzyr08
hHkLm6smcurNJ2WW1ZC8X0pZXSBvNhx2//oYnZvZf9FeobBEbC8eeReTgRR0lnyx
RqFgj1qRhyoT3TIPdzIQnESIlAQn5YU0XoQlrgH87bC5gluoz1qldgq/K3wDbxWd
EDLH+G3cXjClBPL8fbTohVzhPd9HjGXcZ3huge3TmqnLxs/sXwWdlv1O4nWPbFPp
ra1PLC7OsYeeyzv/0swicOqsi7M4mu0JhXnnbtK7Ddnn2fy/7IGLrdphHYy556hH
5Xffc69f7CB0Nyftg/ufHPNh66qoTyHiaTYi9OAScHLMlIbyHk2c0n4FdtA8/4yP
a8Y6nRstNSTA9BRfp7AaIVpe4JON23Hul6P31NGIfz47H5/0+NpINUgJcYhrhEf8
oNwl/dimKrpTPzM/r33y14XS6pY1EelAUM/GUnMqiC+EZ6Vk++L7ZBHmUjj7ED9n
9lPu7D337Yqakbb7IhPsCBzQ5nZzxTkY/zs8JFxFpwUIsYCMXoGV8RrrV1jAtj2y
+WsfQjs9oM1mGjJBx/fp6Sg7emmh1H+ieqOEK3TkMNqmbFHTCDNSbgxPp+hoIxch
sCWbf5l2ZJGJm64BC2x/brbnKW3r5aMEH66vAjGvW76KG/h1jQvs/rpnBFELcswg
IdvlgcRrfJKXaj3YwMRbrCRgnQA1qAt3hb8cXjk/AO3USafEQds+CTSGlbiC/m2h
jdbJpNbBOkZ6S0fsdzaid/VMJr7iP2ZoTpTsLOWH6a1FIanS8BEubljx5hLOwWLI
Bq30KUaYnHAbA1QX0G390kbkUYNyvaCkmXAuv851UDWUSnHziXKMDF4h5OWpbi0M
IC6xKUpXVRvYu3FJFzI0R0WHKJ3KpTVpkIBjPtNeUshKf2cXm2tGw9t/z4Xm/FoT
fX3Hi9WLVG4yIhbeK5/QlJ2Y79zVngo8ejY7TqNG0EOK5iTpja7yEYutJZAwKjD/
WadDoHtnCkc3HlgO20+38t26lao2xpCniqi0ao6e/K+qCljpaZD6DYvzGm60vPJA
o4M6un2OkgPJpTvETRbnVNH0s8iGCkVq0ppvSifygLM3SGRM+eEdvK+oC2sMyxyt
Xu1FAcy9qzZB/48YDzWpoSMr+peeq8AOhw8O6ejHh0nWZ5f1My4ZL11yTJxidgFM
F2lXXXz5Mevj4qdXMvuK9H25+i3ScheKz4FQdVVcfgERzmZHjg9DZPQJpPf3/YSK
2DZYsyWVofMMFcfRtgieT8dQYbhZpJol+wzM75ZxRj38yb/LvZ1uWRu+35XalTRN
sE89SbQUbWFRgsJzjRjwv4ZBiJRW3f2jDEQFd5xJhj0f1UnZJW4f5g35gP/xGKOa
EEHlumtRzsg/RyVYYxD03/hwWvAUV2zIXNhOZCWhloK5lgI43TdjmhG0QW2i+kS9
jxa4DD4k2yw2up4//gv9KSLjPCQRyrCuDCaQVM6EFD7LwbJQTXmW2Y9786nzKFLr
iQ3h+JylxD3RdqSj8Cz3Woqhd3MpIyT1LdXSMCkyH2AUswZrEJSj0QRNiczoL9FT
q6SD307w8bS3EC/Pwt+hRaAu3nHPIFpGDJsTXYjkYzjnU6Ivkew4BF5rtROUOsHZ
+eXo7Emfw4sEO+94zE5sPMQT1KuA7E5SGHzrNxNlDpfSJedK0CbeRVlQ1DnD6Wfo
yhJtE8C9L3p1qGL+VTL4WNHJ4D+/djtIyWNyaqmi40J9Wj3j0aUozudCQY2It/2B
FdFzDVA4RkjZ0JXzGFQcSI6bRoCaPA4Y9wznCf9EJzSLN4sBAAlmJq6vQB5vSqcG
IjxACCuADEWwvgBW6ws3rPJTLUFKdnXdUCAG3Z/4Jw93XysVKcQK07kEsBOgrCDI
QuLSO7Z9BZVxl9dMePqYmGPYx68u90rChGFiLonDBtxcfjR8raQdoW8Oabu0sh7d
sUMU0OIn754pMQQ89mlHkJuuTIX4aLZjHTxiVDqCvZzC2kHXV+LGlOSNE33RPHCT
1w7PEgN4lsimEd7tHdzOCgSBpDp2hsJmVp3Bycj3hoQ9e073Q0Qz5XfLUAGbRdjG
H0pDBD8nbVgEeoKknypZxWp8xzvi42lBUjxIXlt2ZPPF/RbqkPpDaxgWmm7mAKsj
K7So2yJpiOgKmyECNKr4qj2lG8WWGUGGJm1N1RkVidAZJfbabAOqp8YZcAkhY2/q
bI1V76ha/j1LqwJ9yB402x+3HAJ5tvsWS0vrjmqI1XLOOAVE3HBPTGj6/sYl4PK7
MJ+J4jJzzFXobVGrxmed47bCB0Gmmhv2L1nz5chsY9ZSZRJmRv7/mSV57Qp1E0hI
eu7M3uouZgXIcoNlCiKzXJTqN44Rl8xVjmGc5l6cIUDkS1xGZOJeXAMUALlr+7nn
wf0WirGHQz2Z1VqQNV0GwaqxrlHVGOhlQt6oG+4pm4ON7sd/Fwfb9fE5becIqC4y
85NGLkTj1NsnhDjyquzch+a3Ev12FZxyUWSMeL5jQybQXxi928a/6vhXYm87f1Sc
AyyyACcf1YsVXFzC0MfxZYNu/+NNblAgSlg+S8b2tbvQjjIp9gHKm/bsFc2M3neD
DU67sJxROoUY2B2TAOyv9/w3k3E802QJwFscVqPFl7ix79Dug7VdUgre1aPK6ieK
ThqCo7R933cOs3kLlK4B8t3EY7QFodhIxq9D2vTs9txMa2oIwRd5wi4YZPFXifnB
fIpYm63K8krXeGacjC56j5CuT+tI2/XFgVuw6ljnjIDwSr1hKpuytthoBynE+XR0
u0Rs6PodLgrhgBnqPUgSukU70hg94hGPFz1jDrh8aC599qvzx9/dhgDClk6LunK0
8v3tVSiHWl7yyOzu8qNrGtF9HCINiu7IMma5OeDIOqq+1+cQQyT2w+bllvn5Rif4
dyOL5+fPB+VbnUeFAmc70iReEh1mrAoBiK8odsT/oZXi4Ls+2yYBVCerDwzmcR+a
seFJas7bEUkz3oBJ9bNVTAxJvvffpcsUVNQBMViNhm4LoIlZ9bOYqj+BOOAdNTKl
fhaMEkfbgSyu20deuhmdsIcqt5H02MujvpHcKc93kE5VCtx4ipid7uHWMg04ahRV
cFoHS2s9K4cvAn0vmaCukFSkGHcGwuyjL6zFC5YGQPFa2ROrgNsCtQzgPxvQksY2
xTwQsAbL19nuZTjE6j0qtiG33wqjwLGsHGTg6jAu0Sa2PzVZadXo6CZHPJszxu68
Thrf0KhrfFH9pmnptXTHJhhxj0LS+R6uXaagGVmKhEvAqTDXrPsVJ1BHCSd/DGPz
E9zbtSL04JtX7LmC4rnc9NkcSV6mWLtCbzniqA+YpkM2CvkB6oeeJ7GYVi+Ev5ws
J/7B4CDkCB9QlEVCLvtMnK4ZIsO49YPHvE1JflEg4AAV84BQkImPz+Z5b0ZwPJJt
Bp+9ae8CrMDlsRc0ME/7ieJfAi1u2Okjbnb1pRjokHXf5wnCEiqTHVUigDt5eh8R
nNgx6LbxtP9tfq6Ls4RCGv852+z0LqcifbAFbJjmHOsYIx0bpzDGI+wACOiZ7fVJ
anFHUQdcjZq07+wxVJzwkmr3CVyywVLA1CNASkG1+XV5wNgtTXGgI5jFt+WjaMbS
jQ0mTqCMcID9VMqVo2SO537EHHPKEquXmLSUAPXgnhecwpEfyuVUXXIfVD37Nsiq
ec93TCJTgnuknfzPzRGPxLtV7Ae5t9/Mi0U9ljq+ucVtQaNLd6nT+p6kW7UxlUn4
FHuer1bhYq7xt+lotXgFj+K6p52ZpCdSFsl/m5jwtOBhORwFQ1Yovivs71XsweSO
CSaawGaJEl2oiwM2XZoAeJwi98Ehz+P3M85nR6p06si2a6UKoXF9BKu5pY+vGI5I
91c26xUpj2Z42C0BLrTn/vw476VXP7FqhBcS0AHTE0Rcx3V3225mZlZv0Gbi4t0W
QWXe5PsGgeOwxzMXHO5JWtRn7GqpjwlZwacKEbnhKsMKGdDqP5/0Xv9BhWmk9F3r
22Y3MtwwrlVWsGMcKHHr1qjd6mefG/Yu11cbUISrKbxIkqfobxP7KVNFvUOXEP6W
gNENGnC7R7dMljyn3z8NF1H0pJUOWu7H4nWu9q6jJH1JeltvTcrLM8VCgBMz5yMx
BstKrmiDRyDPSohZnE72Rjjn3cAqptAFLjdeUy3RTXWUhaAJ/C4jiQpoGYITRC1A
5Qhl7uUx3MKeI0KASBKxwCofnUhrYwqCLSKpcx7WyzOc3aapFpfmlYN4OHSSFTPx
t6AFKJpaPLw7k8HnwnG+cyZA9CJ2R0m0GOsTAbsEj2ivHcJKwWXleKtbXjIhzPby
WfbAcxXEZ4euGnyqtL9hc3LQ5Cx7twc4MunVaHPKgPQ12pFwwZNFP5zSQoYlvKBE
NOtJ5uibBGqohbHes6tSlhLsaoZoiezSbYJdCiT82CKiVPG2Xtawv/FjXRql4GMT
YgYyaZtPNBTHhsZRgsANfPct6U1dEpqWOaroAz3xCPlgPT0YITU4CSC6slByQliT
upGWc4MtwRqVcGEsxcWrOeyXbbbI6RJ03juuD9K87dbfWZ+bYZiWmVgOPPR5C+Ae
GYXi1ujaodtNwy5vffaLh6yXujoq5+9vzPp9BdtGbbK4S1FobmFcQAm+ZC1W5/xF
zpqDEtQLkd8t3L4rKYG3SDxUeNZcwCifZBMzAdl1p4B+tRFtWWx9Y32zu34mnudc
D5jrRKWdlQhphr1UXUBDjn0meAOdHQblvZbG9JAs2MXrDw9H+h7dkOHa5xwXmPbk
0hiCG6z0mztzotmYMqgCYgDbPte93skkf5FTisyLhD/Ql55euru1XIdA0gBZpq/y
PR6HJcOgP9JItNhASti+UdaKR+JOqDCpEvv7NpYMy5h2IlVIoTxwgWwEHC+huKxO
+jKgfSQqAOKF2+ZDVPK9r3C6/VbZ21RunGBIcJyj3/AAvWaj+hO9LFNi2SQzs7vn
XI0eyHUuOIqXPzJhvHHMOwU6YsO/jOGPruCW9S/sCT7jFp20KSNJXETKQNO3y/+s
FcpldvFcpk6kyW0x/nD2mmXZx+AWLZ6pHDw/YqLTyfisYtzprzwoi0M3C3pTj0Wy
qZJVGQ+t9L3UBRhBMdlv+BGR3nv+il12ntXbsOPbYSK8ktXKNtUhPb3iFkvp78ZQ
/T83dPWWPSL98qW/suR9i62ZElPn8GZ8NpkAfBBMmtdL3MuDg+4F3EfTlhUhFM3u
MO2/pCbNR5Yv6rt961j0Lj/f/OCh+r3LSW0BDDul4NUxaUa1Gw2F6l3KwmXteWaf
Ri2a2cwank1QK+hwGx9v2K/2Rdl4AjMwzzYDV6UAJuu9TbM15cWZtUi3xo1RUuiq
NFPNOK4VliobfD6EWbkDW+SJbHvsmBa/6QpuB7qeELnCAKMlqYXILmMPl82/KYtD
kY1AcQCKEg2FJqh47S370+OVO8FQbRQ5c8rONMMbw6SweCEUMP6NYwBtDCKHaVB8
PKFrldOZ4M0eJMk1r1wq8RQOtMomWiQOqcdzoli3y7T3XiBoFHprHqm6eyy1ZxqO
wj/vkq/qI99ORfiOCr8nYMKucgRfmkS1w2bjxJeliA5RZOxmjFTEGJfZT/sebAtF
FsWvUW8u1wqMUbANonPHD3ptgtDvoUDsG7kEwrCeH7jy8WyUczucRBFuBbS0GJth
uTNUvPTme67fSEVm7zsaGVeWCzHDkm44TS5W6heR8txXGM9ap1yqoD09mVII/wSG
AEhjIMhUV2wce897EM8sH98eiRxFDWCjGuQ/IVzBdWTef+ATQVF5ZgkeV9dah2fs
ZmARxqNKOz+I6bPKlFh4rlewQi7M7jrWWuz3MKnK8qWoeHcoKG4cazkHrACaXVTZ
99Rgnksh1ZfDis0OoE378fF4caDu1aML5CjXvI8D6CHNwYEcCZyabveRVyWXyVrT
FC0s7VMlgl4150hKMa7xoVxffr4S7yW71+gUM63csy0nY30s8MSzDSgDxFMcHsre
9yTBXfI0cX8EV5yt6j7v3pjnsZP4fgTo97SmJFfvAK+ugE+dEYoEwvuAea9tgjdo
UiLSfqW1UeYPDtQ/QLzl+2nrxXc0FVr4DcqxR2fYzyt9+v8yD8INYpw36+3OGtH2
SdaHMvrukitOCydWZvft3mw1Q816RObwu2qGIgnowDlkvmmtqZZwTZ3LvU/auylf
3xKMJxWLOaWOvfWbOq7PbiH7B5L3bqkc9D4YUVTo7I+dzbBZRYY10zrG0eHy6bkd
toO99Vkf+YvI1lHaqV+Rl0S7BVv2x8XGN7x6z+7t7xhk41oNJumOJNanhkcEDQAz
gceYasVH4hKirWaFqkKl09TaMekMt2qcK8TmqUCjkQYHE444vyRTcz6oXCuSwIwS
YZHKIrikQDJHfPAodQmFmbwG7+7emSIGKcdswG2Euyme41WFNJfVSaaIlVLtypuc
cAJGeUHoSrQxoyXtFeghY4VVE31tjPHaJviJwG8HGbJ6MupyehV9OebWOR6Iban6
es4zwzRNUSd4gaM4nwx1FS9LYz078Ncf8oNXgOg7Y9z65Bni30Arol2/Hu8CqnXl
nKEeK+M1716OQUXWZ+Cv2NrtCdppX72ddS1mzUiCuK3eUpoLGu/W5bYd0vQsEDGe
njtThRaPtSDwjxoi2rD7wtyyEj62JZT+0yXKmScRcwIo4ThXB3TUUDApDweafRpr
d3idz+6vl69WP9ThDZr99/ZYgNA6UMUnd79FETwOMDOV9GJDBMw26rzbzZz9zBSK
ZGxMYDtJZVYsGj6FaS4bQBPjUJQyEgtheNAu2qvNzDgKDU5prn64awbR66XjuqH1
I0ZLsh/GP66TBb32ZLQf9hdlTnfHVhh3nbKM2Oq1hdKnwvUc77NLQWRaawz0+Dit
typa7sw8Y8Oqr3KMkLysD6ac8DZCTDKGLQrlB/4f+NPGAbpltGvO6QgfTWxRkur8
GaI6kEEQiwgUAq7bSrJvAwijeqMTxnwqFmXvvU3lECnJTIKnS7n3HnG78YJp8h6e
s2q9o2h3+Ff53BOxvPDk16GurxAPma7XwDthK5BPfbYpn9Lr5Bhvre4GjOo9qVsq
esRb97+ibQDF4PBCzYYV3BExEn0J+5TjEpDasfGezCU+LC9BUbH19vMChqkMvyRK
LpVo3xndXCltkhWvDX8Zcyq4dAz6ZSpn++2LQBk+HVDvTQvkZgmK/iH1mPtgtHLr
I1MAiJ5UV5NJ0yx1HO1414FPBG9GnZs8qZVlu8ZVyYTLh3SCZUFmsLeCTf35Hi7U
yXU09zs+IH1KNde1ib7b37iwrsCtYgYXY1jiTgzhsZwDPVm/ofpw/tL+ox0cnMAs
D0ZM0gbceEA+zvo2iTWhyPK5ZEw6mOrWbvFg/TSglus6yh6PG4EBSHCQZ2IjcmIF
RSwJyjgwMVFD1NpdxSUEotbdGuqcYGp24ci0kLqrCSpSSuxt3XpcQb4xQ95Xux1m
x2ExtHLY/LsftbkIKd/5ZK+Lt56TwIHzUXgd4Lx81bNASf1yPJGQlUp9UkIoQIIZ
I1KS17iXFh+6ii8UZfKJzLsODR9zuLExl70j8XzqXXYbqwfvQiB8iAW9VXAcoKzV
LU+chgYJZJqwlGAOpWtKCJu6reXM4ARgPGkBRTsUMM7wtN2BeHlkX3MqcNMCUMSW
OQRNrQRIBtsGZbxvD633TIIwU0fyKCmwiEf1ixpD+uhLGY+oxRiqym2actSt9Ea7
FJnzZl9kNG+40Ho2NASF8Ftx/Qw2BgjWSE5sfJSDjFRAHzRuUHlV4iKFukkL3RJM
Q94EgUFpr9UOjOQhLX1mOQm+BRf87qxd0vrCE2HX/HutggFn4oBr5w2crYtTy/KN
jDEgHN5WsZMIQ7OOVVLmfpIwabv8CO42Uk5L4QAUd5pzVZjhQ9vvFEHt5RK2oPah
+pdxGrLblm69o2GnaeVl6tKO/us3DtNuor0XetDfewxDphjPuH+O+bYe+InZVhb9
s802Um5zJbivk5ex9V4bAHIzZPyClXRcXG2KmOvG6DHxGf8TYPFdfob8NyyrGHpl
DVgqpOw5DplZAKVjhqn6lBD8wRTBUXf3adSXjDIzqJ/2SikF2pup40F14MfBpp3f
WA3iDnW3J/FSNv6uVfQ01ztuZIQh8Lihp9Ge0gEDPtCFUwvSCeUGIeG56z+1DoI7
FrvZbqRukLgHpjvqSpS82+Rq9P3FFQ4FjtajCibErVYQox4S6AtOsOaarYYvpCW/
bKweMjdrmojVd+DKQZdbUqoa8EDBYLTveJm1B06ExUSIzU8w1ph3Tn7PMcfH90s0
xjMi/09xNFwyj+u1rxN3zOcRy0DSSSkexYmqcF1+X8g3/HS0qaEpqxGZBkfskq8L
Zmwd0+peM1Q8hHxakw8ZeVR8wuB7BvWZd1E+Vlmfjvt8Aqt1Jf8M0+MWpk4XbJny
EXLl1QCENXBy0rpZxD3rCnAmbX06EzwJSqggxUU28cZWMqOODO8d2drMP5nxmLSm
wxAnOqKmJmGlg3vc6LwiS0P6cC5nsAD1iXcvSnwVsX39F5tUdKGsr/GEOa99M6xK
+TWQxIIPOL43v2sCEonwOxw+z9dh/1OIBpGpZnQR/w8=
`protect END_PROTECTED
