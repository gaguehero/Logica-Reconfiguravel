`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gLQnuFCUuY1oiP6vP99WSqHj0e1cnjjMK0Sh0E5YW2zV9BRJwYlg3gAMbn/Y1us
+hoXY6Yy+vMAu+aH0CjC1jnDhGg+CH9lGhIQJBLSsm50NajR/63TVMQ+NYZ6CZgm
dhw8mW7R+ypXwJlb6EOvaWjpOmryw0JAatRhsamsaDmaJ+eIbEEojXoTPGyhdhz/
UInkF0cmPsvuoIequmbU5l9e5Pe6LVG4NxAqwkbybuReH71vzlbDj8Re5o81pgnU
EcRCzuMH2gS99DM5QMwFTjsbRr89kkdSl7Sbg0/GPIkRKiU4yf96RrY99iIkry48
5TfcLfaPSxeEPZ5T4ZOu0S0dTsHfkR7NByeiwZ/gQbXNDlDfEJ1qwxsI8d8iplAW
e3Hw2ltDrLv+vXNNYNeM+p4UNgfDcVwdG/ahZJ22r7IB3zAvrletaGNOK3OevCcs
qYjsnqw1wwSnpwUXR0SwoVolo6VELiuni88n/fzgv9GZOreRQWmr1R8/nPVrPRfk
yDJlCRfGxnCec2ttqRFHnvaaZWg3VCF8FDhuZwexEq+4vR3r3CJwysI8aqfJygqn
v1MzAXXpgeVnpvdrCQMqAv/lhTaWdH902ztoMrhxnIhOQhQmoKNw4093q4W4jweR
CNOKcG6SMmdMONaamHSYeVk4rO+hxoAZ4wfbtmGcpT8QEO2xkMjkCZTv8562q8oZ
e1yaDrFyKX/LtqepJ/KBv8bZd6tnw9PPYSZuFWbpAGNsChPCs1HqE093cENx4shi
Jo9YpiC/sbM7f3uMEbSjJLCEe5GXaPqQUVtxXNpAoGurhCXHpjli+joGDd3+im3W
3sU9oTjNbp72+xANkWom4vRA4svtFAWctk2yHC3tSnPnrp4+cBuOcfN6WMb8e2Wl
dJcdTmAf3N77RiMJjhZWECb6qhI3ms5Tf3dsNX1pGoK5vdoH+BiZE8TQHdoRAmOZ
phF+H/1h9JhLmVovBjkNe6bCIm8Y5kImD4JOUkUiaPm82pr8j5lydYk3gljb8tLD
ndxdwJPVkwnI9he9rWYknl/m/zChbJO4ZBy9lJV+iAHWg7JMCBo1hIQ2U/Fynfrx
TdtQ1gpuc5rrF6pvez0KNCx6yYKKCd5F5BJG3adsn4nBW24QOUedC6w6X9nTTxPN
usEqhKEJXy6kVhwjh8fqDHh476nT68wWIeiYy4V1NbJ1nEAbYUq4ZR2daJ2OdDf0
raP7b5lo06zdC38+9OSoNIIkM4ZxIFJVjEgBta3Z9JQl8eMmAYd7+R2u2aUncGkb
qiT9uedQ8g312P6aUfkhoLmgxH1Yl06WHKA0yrb2onA/dFF1pfekC4WAamAKAVbY
mPsdv1P9kVUToTUHwJbX8fbUtXf8QhKr7OnQAWoXHElL7WDV6bIssNXUQw2NGSVy
4sWrraaqoa6iiue+mXXn1tTLEvQwJ1TxMEpcDoZWiS6VmCdBDfDokCo3K5hz58Rv
AVcZFg8OjKCYmU1NiXphUe3sDMzX9jfPjFUbUg7VuM4aaNci5HoK8D6C2iY7cYsK
8cuz5JW0HNRwZIEwqE6MhKx51FwzyvzVby+MqdlsvfDWqsLZpEkSIurdCX280LC8
j/lJG6nhcBe2Dm1FArShyuZIjMH6V7PEYYFJrm0B/nscnCpXYIKzi/LQDbedjM4V
amRFK6osHGSqGCTBb3e+38TxvlF5UHfqsDbPvNHtjE3PidTkCj1UWJ8Tx7HvqStX
axL5HE6kOB5xQl5FzmxSssYVf1XpZ0T5kMKY9ktjy3/zul2KTDNydTDfk3TUuMVJ
cmSQEB8AveHVkl08bBc8qcq5WjXGQj4fLvwMUYQNTagQqTDRPvcLFsxeaaXxAs3Q
QBLKYphIEqSF1log3EfmGgay0F8qGGm3EwpwyZdWtFvZAJ25+a4qLCYEM7LCpjcx
U8kt/eKFHYs1OrYidoahCYy2Pq2vYOMoXMm+QqDwhwxj2jlxy24HMnDTpTCeL/95
eDeM/wPK9gqdD7pMAJiWcg==
`protect END_PROTECTED
