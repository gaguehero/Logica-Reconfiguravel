`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yM5NJ5NbKug8eYQEf/qYLrEx0MgqV+PzOhOhssdz+uv9BdgBEcmw47W5x7GbSH+a
Dl90WJgQLd6EI0lG/4+euP8odeGV2qqpBJY6gqAASVSP64A6jJtQj3eLssUBukqW
2JMrDLJVLMEbc80fGiG+yLCKMNlL4fZM0aPYKbrBRb/moeE6p545/ZH5VZULQ5DD
qQaduKzoI8EexGR5/1r7ET0VGBNJY1uk9C46ynK88FQ5YIYrC90UzbAc3dMtTXVn
nMa0CjSRbuwZv3ehpSwB2wXne1HNM2EcUuea+C90bvtkKBQi8acP8P4XkpcI2Q0Z
7UDviy07gHZEeeXqciQ9O76M89BA0FucnPFFrP2xvfwXPDroy46/AfHkNm0vxxkj
lYQupl79GeJNUZRRkMjZO7N+Drfhlk2CpMag8HT38JkdmUEKkblPPWFsYeJkyhvd
8q5BILMGLZHbqXSJCXsgnOKAA3kiruFVQLjbt2dR4D1o1te/mUw9oAtaeUecUzRh
XxGUAuvh1rAeOaKD37UPyWnDaSpgKkkiAV2HdL8z/ffeBo9Jl6k2Yir4dO5uJn0V
o0DXCTn/Sf40AQ7zjgwktn1KG+KvqiJQsEYxSvqjNNPxiKwYfwYkK6FuGPc45U1t
l+n1jdD54HTFh1j3iai/a/+4WOJ65Xg3E0lz8xQYGrKpCPzyxE9RoUrUPmHwwtrB
D7NNMUkb0vo2RurWJbYYGtn1vDsSl0Vlpw1Z+GMKxRElg7IkRkG/OOL6laaU0eHu
vc+t5cN2YH+ViySeyFCkqXjNZ2C8BwgVMsJP2Hccr90Y2KDQGceO5aRh+oqICG9C
s52laVy4PNob1MZ4asWhBychJBDVAvlFdbLYjTyCBThDcqmp0Zj55PULYSxXPa9V
qtISRWiduGm4/p77cz2bsPhfqa+mz87616ZmQzvd2VZ3LGX3vP28qTlRtu9K2pBc
kj9E3jNiJw7LLcaFSQXEytik8pq9N7v/jl7Q0ak/s6TcL7dVDp1hMDJqLjMvWnDO
s7aq8i0ynSU+1JbJIAHB1BeyrFVV1OLhzJvOdFyabY1OORK6Ayj+aJslsZsXuXrR
5IN8pjjpAzNPwQPzYfHpuXNcnQeGkqzBYDM47VLu607EMyZQfTP+c0GQZrNG6n1E
CHTEap1Yx2PJ5Jjiz0S2feGNRoIWH3Kfy1KxwXh1Mno2lvmPt2kPIPV6IKJDsBdD
XHk/CiuV3Frh8fVkHl+6pCOKKkvZpOuf//nixY7mjFdTtiBhLGs30W2hLpryqVXl
LJX4sqPVxO/KtopDb9zNTybcWJdts6bZR8w0dA6p/hMOmyxtwqnqChYzC70dJbBc
69BH/trCpRJytumgBIDEPhesXV0ZXIdIY3H4/MHZHmwLVJU5Ttoqs+vvcfGAd1pX
KYzvK0eg9zD4QesWT1+WdFvKVuHoa4ILVYbuiJWUJE+xomLuQojUE2DRyRIpHNEk
trBycFq8jTGBKhQFO7LJ9CBWclD7u7Eb+CnwCMZ3FDVMP+c/RXebNlXoSEurKGgb
TcMT2LHFcDtKLPj9LwAS1Kokk83NPVpMavl9gZBrIjT4Bl3z/RZI4+TQM5malmeu
J5QkG+PyKh6wL3zJ8j2v9nyMdGwbMRzcyuOqT+cWmT0AabRd3afsI9PetVQ8MYA3
FvnpNV5M66EyGJGaZY7vw4T2SFYPe427TVu42s+YIW17JTXlM3IPHh5TSzlmIh8Q
yGFC9lSOT8DG4FMxB8xs0PvlXO3rs97JS+/Qvo7mBd5Vdj4bZT63KUZ48Sew8VaT
G8cRXIgFpa+3K+elgcxXMRGfXlEn55v4CBJOnUQtgVYNuKdtq1AoygSBEw1RqHTj
BVoTuLHZ1YQLyJcCpqerrfmwNozb89EzFnWEpIY80iQwIgHqdW4f1dO3Q8G413CS
KOtGBuwYq8slCMK/8E39kNnhh4qmbn9apbUYNrUBpGy8LQ85vQYZJi08p8s3hP1C
7bWreCiqzDe/bccc7bLgZAusowHiIItclJ1WpJlwX0LkQ6lYMfgCTSq54MWr/dMw
`protect END_PROTECTED
