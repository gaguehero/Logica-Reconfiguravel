`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ioTGKe2FX02W3+x4YoDjS2gQxutYnkM5q1e4ybYDPIFvPseqsyBePXxb6tDY+9bi
62VXoCrbh5l+OMS74/IjVn2Gv62EumLS083O24McGt4D6HOybGv+4Oe+OEItV1kY
QJD6CMpj69ZHexlHL+uZu5Lksvu94rxEvxZX009X2pX9Na7RpUzhlc2Se8pUBwN9
f3t28y+lSZZXg2mJNH6vXiBcq4QQKtGgVWGteDd5a7QVml3VolLD3Tl+rgUHZy5f
gqifmmlfEEzGPWlRhvFDhcgSMsiq2X8jdvvvLVyRlFCNdASXW+WmpFr0oCE9cZU9
v86euAm4gcirkHW+eC/tH4OMQQfXTQbIxwZX98DhVOqfM1ExRMyjVaqZMHjKai2v
PpTkjQpuJDxe3p6rW2amlVslwqtEVqqBHmjhPbBqHJId2RzEtaBazdIP9vDZwQUp
yner7SN1ywoFWgzMHc2jf2TdS6MWubJtBrSu08jSjjI5fGDB2m0trOhWMF/pykW4
FE2aJT471SI+TdQRN7RaSc3msvaWnTBitw8hQP93us3m5rlwYuoEo8x06V9+rOKy
sYBE5Cn9XrVcuPc+ZYZifxj0qtLBeW+aqQ/zQbBaQS2Gv3YV8cD50xsBRUxs+JvA
PcpAjQVNmX1AbQyHfWnOSPqPO+TE6D2Ba0lC31OAcH81bG94cjugd/f80FCPq6UK
Y6stUJqPEjvPpKtai6dR11Us6Mb6a9Y9JmsKD9TnzMUOCGnshQ5KdUNPenJzlXpC
ji/mXl3Jbqh5dHEEkilzDNf9fhXcNRzLQVmDw+q6Ev7AnPcGDICxQPLLj+axE5Zc
zB2TkkJZg+NI0y9Ci62Fkub3dBrZ0FURIDYVUsttZpkWJ3eK3cSeaocHSymj5Ejt
9qASQy9jkdnF7YAXyt0lNqGDO1MQqXX2JD7FPhEuJyVNEoet2N3ohUGFDpfuYfwt
vhCGtxV3oM+Ii6Xp2PpJ19C8UCnYr5eWiT3573phXaInDiROfzuNk5+3EflkiieO
wziQzQEKFASlHZnkG0hmvYC/qZEw2nxF9u6Zr7mw0S+16U9wunVTgHgNVbPLXRYr
yHwd4MSkFtaWxsf8f9EDHovSq5S0Hp7PMAbbwuc4V4PbcUD2tJoi77IASm1cak3g
NVjlBMoPHBYK6lvWLjxhvEWSQHDvdESx/m9O2m7cx1c9TtRaAPHAOZLIujH8j8Ln
dqGNG2Ki1VMaaAsO0oXFlQfSqmts2rDeMdeU+8JF6xNd5fYbLzlQKK/GgZLUcCGj
ZRhX8hr0mdOMWATtHODQEp5HMqeyNNJ8DKtX481Dwq4sK+xj3Op/50irvRLA/2z3
p5A9XZd7Rm6L5e3HRXpkkWGB/0JfoT4/xftB5+x5vSaKdratzaw+LYYJO8h04Eck
6prL7vILYXIawiDxyLQ0EeqwM2ExPmpfVuPL9jTe1tubvPwSdo5RELSi8wEWUSM+
nNHxwJ6LKH9AuGd9XonPh/3H82W8+YHqx9chXMyPwcGOyLK3ARqDtje+WVE/8IS9
kf6gmgdy1PWoib8nADcvd/J9JjQg81MvjqPVv5bLkUrZPxhmM2OzCvednBVzxdg4
nOYhwS60NK+b5ul7R/CD1BdBx4P71+4mnIU1SFQfnGNXFgg4jN0sgd39j4cb46Fb
QvjoVPeFs1CLDmWn91G2Myz6TWNXR6RKNRTRCYHf34vOZTJnwmf2gEveI69rIfcS
loU8P3At4QliAIvtwhkaIpe43bN7TmoSrjWpDixXcARaovFPmPBjHvJHpzkdOvgz
gnVREECUrWx4mOg7u0E62G/SKuVnniAL2eB0eLgxQmP+PlR8DXfdqgFPpIV7W8l1
PAqmwtHV4YquoDsB/HN15TKr/hTYMnVPNCAXLlV2qI0aawd0zXNGhvMtcRWkiHo2
2k0pz2SIVyt+1Il3o3Xya4dMBXVOxu9I9tbUFKpdhN0oYSbUxh7kinNBoAB6ROtn
80pbr/tRuOxRHtNjWkczKIHQe4bxlTwXykv/2vdGzHQqrWaFlqJMyPMBYKmnGN4I
qtZZwGbcY8/V79BnNH8rPJ18tJulpKfDcIYyEoLh6TzyTxVl5hH7SL/B3p2mnvbX
ppnV2+Sd+kb/JI1rlUqLVaruBU5eFuwTZAc++xOcugtgAXiSLRGzurfREX1mjXSk
vGBD5jhdj/bjc0iNlzAWPS8ezfw1XW2AyzbZlQks0fxKFL5ISQtXKNPdYFENXUk5
IwsuhLvUDY1WZjkwuLiIEq8ExonqP9dxhHc+ABvygoPiUcq+e9pU6VXXom0JIyYm
JXYrrNqYqQvNJW284xo09vD0baNs6hwrGb9g/LafoUf8ipe2Pa7Ygg3oNgmfJT0S
tg/SDGVoppM3e9sxYzldh498Yn49k9RzcyIMPFxQ+WTQoG92ljhJdjH92/OC1Vkj
ucKbI5Ga5h/BjW0A/n6bcYBAaYmEo3HxFNksaqCzdCYC8KEnXMW3F9xfuHaWtizM
myT4ShepbHwbTm06x7tM2fsbKYA+EXaCtutfJd3/RWh/vluZrai3/0dvFINYK740
oo0weMDsWXF35WbAvAvzxIs97pVVQMyhVGHRKQSKjaARhjYISylskvGIiO0rOdQU
LfZityG3pVKr6iKX43GFXWhDc0IhlAz+QhSL4/DbIputlQtXRKUZMXlOzjE3iLn6
pP9Av3DnNsgEVqY9VKbdqac4KU4vM4F4sG7ayydbLpJc8RB3hmPNIbqe9i9GcVV4
urZNXfUjsIf8c+1NfToPxMG+k/VO2oi2ZmtKn3gKuyYBmrtyr/JPl13ZixeemPn8
UnJngPbCkhJ6dzAviRZUP9qj1uc0DPDnkGkw6fVFrE3mjpo2kcsIrQvquZulzIji
N6DeXs0TPc7L1sUncO+kO9eiz2ol5TKIEb5JB0w8/SU3sh67zhZ0SKp94HNMZ6W/
MHQe+RK5cwZPpWda3AphhRYFKC4c+AfcXmXziyXfhEeNc/QM7AvAy4wu0rl5AlEn
xOUM3GYsN6t268/KXaOmWyPq/SULKLFtwdXnAtNmNXqlGbc37IPj65PtSmnfGob4
O+9eblIB7hFiD+wFQUa7nU9+Ad4IGejpgKkY3AWdgD/fmvvsCp/6EgxI2BkyxZN+
WQ47bI10GuMI3Cl/LYvEuOf9YDPEC+4RbxTMsVGKb3x46IPL7cTDHPMayHdkwnUs
detKxwJckdsqmav6QTp2eQ6C8PJvkJQay10EpATC5qHJogJ5Psy5DRT4CbJcaFfy
Odtv7tA9kt3kj7MqU09WqRMdLub4fg36GPIrYTXVNE4PQaI2zdzZaYz1TgaRGnZz
gXY39LyNydjnz9GxuUN/RRkcPCm3+GcY8PRoCMMkb4D7FERuNyAzhDtnnMkvhg7Y
Huc9HG2FQf7pCfw1dwN6CBwqP0ILr9gRIk3htVgS7M+XSHEeycr2tweT8LyV6AtY
X9QA9cJgWRWDnkyRtKsspcwoMwNN5VU2AycKYbVsSCpWG5Lz9p+DSg88PDcyDITs
itxzE0pgS9fhoi0G5Ry/Vj6avh1GC8fsfJw8tyGbDuQJFiQfGfHmHr8yeKjkjfyM
0pegkVSZarV0LIH8HW8Umh/Oj2VZk7NAIXFXbIK0Tkxfs/dl9SAFLFd/jot8xN8p
M1pVpGP63c2nEBrOsi1CFQVsaem/WHBbGnG81dsuPboCUYPyTygkM8dJffgxso/y
vxZCSB5CkmcxkJ3Ux7AUTB/k998o+HSndAtj9TZU3hbLoTJML2XpwuTG5ais0jJO
QJV/ZCwTkIs8jPw+wxJYTcPO3gufMaqviK5Q7FkK8bFoaLC7PuyzDc/6po0tjto1
rJjX0b8FeSI1HalNzu2i74DM/YNdQO3cpcm20LMJ2WzGbFHP3ggU8xxaEVoTkUNX
hH6u/QmJYs52E4wjGlDIuQafg/AaDSnIVcuZCDxKBM4huWl8IfdruauzH5q7/QSP
tAHZXDC76wsFNyrGQ9EQEtSxbj7dQ3k9WzMCnEvsrxqMRq20yrv3WRyYOqMw+JxY
UTT4ud10T8v/te/h/tfuYkU6Tn7WF5N5HirtA2jsbaFC9070hPPb8M58hpY1EFNV
pyTCjdeprJ2H6VW0NZ1FbTX/iziLUI6t0D0HdSwuZ3qByDEe9nB/ybaj5QicF3dK
+/tVRCYcbxS8SQ08DRwFGDGCX1YDb9qd2AXqrrlXGpwBwruJLKi5jywh/W8PXDSR
Odayvm8uH0pFXdShCw4/+U7wNbpO2+WHj55ElFlgLsGRO+oeNbQBsFXB9k+oPs5B
Ho89LHytvHb4Q6EK1dDcai4ADfHBRdASvaKq5DsF20L592wYXDEU3oTVdNdXHuhq
n654h+G0X5R5PlytQHyqCznEOVbgjKJ2a5YlHjF/OUmgRLGLuSEtF3XU3oV4bgJ7
apsdz2mSAGg6MEC3WtrzSicC5QCRMEaHOAGFr8ooaiEiGdHVmMofS5BEhOlOlWuH
wVYvlbH9lWAQkn1iDAC7+CtypRVwLuPFxLh/2M9bOLLpSiB0EF8156tgb/EL7rDS
rFhC9WA9j5sHHGOVWKCpufqXvC16Gp1AxFzJ6455TBpEMX3G1a0C/Jp0o0iZECrX
opy2QBPkyhoAWFJgfGm8w1oHNGdhqX0Joacn4kBXiLkZgGa0T6N2QteWBEw/I5vG
bIkeJKOYXXsq9c7OuPQlsmUFAMIXiM80CEyKqZinEkL6d8SUuV9/pdXqTpHIbNZY
nWy1DMB01JqwpV4FaZr6IIhsMDoXyJ8TE++QIh1f1VYwEQkoCcXr8L1hD+WLl+3R
8XRs3k0cbycONzU4BxaU3FjDsJDJEbmcL28xubp1XIcHDqeaHUVOumyGBEadM79t
+42+Xz/fgebWrOEZcY/1n3FVPPEVPUAk3+OaYvPlFYIapIDwWP1azOyp0aTxoOJ4
1iosVE1s3b41FO3I0t8I1tFR5v3LBh1XTbBHXYbXL5GiXFfE9TlGkB1xMtlj6p2O
+sfC1mUIyPtP9ubcq2Bv+7n02DmXnutHHfVke7eQnKbqvnjswB3xFB/NWK1oss7F
pwsOf7IPa1WbhnIzx1Qt5JLc8Buj89BLURzwlAS+/43bGMNWMule65Ja8DRlZxc6
PoHB/d7gcn6lAxG+2hp1DgXvTkX+iyNI1nb8eTCQoPa26XFGTouRQ59WRDSib+9l
FWdBCczAJqX3HqpjG7xpp/Dm+xwN5j7fRIY/j/pqYvMIlBdBYNQqGFUq+BjYWJkf
G2S/a4CPQembn6TTY0KBgLp1NAYwSUttV2q6TlcB3wVmANIhzsPuIq2WhuvmMatH
bS93AjVN47k1RKyPORja45aLmp2u70BzYCX6s50gBFqQ+jgVc1wVy+3LiStHQmCr
mAds2tnYen6g6CugiC0E0jkq1qkcTf/fKTbPYOhBlLJsZIVIFI3YXi+4YSDkZ6t4
QNEAGgkeSX/R3Dyuy5WhEfHY0EKAf3uNqXcgFE0WnmDWdrfPBiPHHQLjG6C2NdIo
6OextMp7DxI6vajCQeG5Ja3Pu0GuAdLroaylkl8CWrKgnJNRJ5ypHC5oNiLA1s7Z
ZPWx6emoJtyFcOljJLq9Ii4xXEo6w6+IISi5o60lP/vP/MlSjNPsd30RPUMRJ0RJ
jNOfqHYbAR+BKtoTOoHUxMoD1G9Se65x6UbwPKsrIbQwcD7cvqde/psWDyfI7IPR
MS19ax+BX1mphMU6QIojXmYwVHsVBShGHTjuRn4TTLsFWHKw2yX+piZZMJx/XvwK
pJ5F9WL3cwuY36YuRy0kfqtN12VHUK0GJVaWgzx5va86pSqSGkgnRtq0dEnMXa5w
m1KjAVxLew25Yb9IjAFcXTxMuANveb3BWu7VfE0MY/N9j3eKoWiuRYA+SN73xQJQ
wWTFU00/NwE7lklSdoDMgw2fbSMlgyt50FP6tcDpnU/jilnm37wBGStQYSmPfnd3
DMmGQYKJRJOGTcE+uPnFX8quwI/CmeO2tPldTfFckvuOLzYjIBsNp70YkmXTOz1V
zDeSUmWnsvcjw05BZxySc2ywFMzvh6YSNkcle11tslMKienho3S3uYiS7Pqg5LQc
1kZSxRBAn+aUbq0ns4qyc2LDaZQPqWBEM7xmYAbgPF+mli8F2JGDriJa1rKumIYB
NYpUDC9b4xuIQnW6XfC7vPcNxzuGlVFfA6RQmw79UGJxmEPDIbcojkEuKcVim9Gi
onX+xbnU1EqlFrpVozpnjGyrVE0exOK3UtEfjSRmMNTpMMLQtP5N4t72YiJsEpns
sEo9VPEslRFOxIbO7Q47dXAhCMdr9HKGNOGhIfcxhPsioEVW/j8G51x/aWvMhwol
3nhVVKp6MWlpsudnTKYtMYLlzoVmrwk5fdbZQKVnnNvWu4eqWxtvJOOcufIn6Jun
FM/tqx0nEEE9I9AQZ9EDLlzqtDNX/ESyBMwtnqI2FwJ/OZ4ku4VvjRT1FYNW9BSZ
r2PlvUDlR4PhLsC8TAMto1hfVvY2Kd5s5VU0CggXmc7qhAFD2nxuK5S4T/p7BCGx
hpamAY/hvpy6UwAlT04IOSMxDgu7rWpv4NwH1haqSCeAGdW5fIVqkwvTiozhzLTJ
asUaApDNfBKdeQOU7gsEPFmlnQqZ8m269s2w8SRXqnWNyMz5BbrNVGOlZfAZzP8a
YZaIGl6FiOPTOVRqaNnIVTjgqU5YH5t0Fd3sA6D1Yk5AASuv+3HiYTh1/zmVZHTo
YASEKdBocnemGISF8bdw7Y5eieECdXc0banHZ31Rk72/ycvBJ4/1XZT0TPFfdkRQ
X5uu08gyc1ubx4jVfL6/s4bsYf2xtU6nvaTS6ViofaoGooclSHBoOlw6BxvxQ4/O
RhHbo2/iYS1tukpOxhYPGu/I1BzBO3ndXzciTIQjVzYv5vX21X/P3bM2QQLVpxoX
F0rLZG6ZdR0Fzc10YQs5E0jhXeZcWXFRsO+IdNfNZjYXA7rR+bUeTucEc1PecaGw
LI0KqQNsr0Ev6fw6zgfjqBTgEytCW+x1oLUk4ZsZUjLpF3a3Fmr5/uw7iWQoWTaG
CKE9h2twTkQwifEh6kQ9g3IfCZ+BQrf8kFXudh4TYHVeudRacm7lsHwGvvC2NI3x
B0hi/mB/zDPeo7LWnjKLJcmSsX1TKt9BOSbHvJAlBHW+GTzuLvFHRgC8OhJpYk+f
r+tkCMgOA/ECgGQh1sIHkR5ON23h4i5k7xUxFrmXkISmCpmeZ1NATcC8DhENfROc
lp5MHMudlf9hY1vSbq+tnIT0GySxBnsaUF7bhGkz0zUXumKA8XkEwvZxGazuVjbb
kGtZ+YhRg3RNVRaw0wCcSMi/Qq73puFVq0wvg/p+UGCPpZOE+kV3+OP24Grrnp0e
Q8v78kE92ZbLt++hDEdqxKt1u/2fBhVcovR28f3OoJTjqA8ha9i8HwYBaOKDvnMJ
N9eFUVyke9Ns462N21cX+sqgDtju5OwBxMYxuLYUlSsjh/nu+j6W13xn8P6qGjtl
0sxXu7zbiONlS84/jYkfQoywYUTY3k2KwHp/CzI+tjURW8E1enfYghmB85nn1Pe0
brRTvf+p36zTP9HXnV/ItkexqAp57gjM8MDAVmxI5sG+SiAGZzvOB7saGzfr1Y5h
8nBz680ud6LrrGT5SXawe22CH1pZAHAa1CHvYRxEt9I2YuSXBu4FVT3xW45mfWuQ
`protect END_PROTECTED
