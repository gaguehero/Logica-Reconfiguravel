`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWqW65txpku4vesVykcUP7mfM41He/apMQNLIzeobP0UUYV4U9DJNGoe2Sx8oDr4
2H1eZULQAu43howQwdyEKdwZAdapHO5iwpCF1mtzfAENgPUsjbPN7yu8Gg+xurHD
CaceD2GxDReW3Z4d+QPGeUj2sgb2y5e6KZAqpEierNE4gnQaxL9OVIM8LDSRmUjs
IjH7C6DX9AVO49vtM6n6+g/9YpQpE5JlwnNgaVQswOrvCYYocrwgwU2FB4M+TGul
+pKXeN2q1hFIIg2djSaWElnVXaDkgASvhM+osLy8dT5fv19GGld/QDv1mm49G5yO
naP6KVxdxaPIMA4Nl9f+l+QHXMfdY/zAuftukg8DJyjW/l3yTnbPLNCOXnDklFu9
s2QQLurCjrSJsvu3QSA5B9C/m00/oSLDZf/pWOoNjAudX6zJaOvnDA0d1aeS1NCC
czmYhPfKwpYmoeC5Y8U/kiHHaLYZrUqScrATD3KN5/UPYHuliKVxdLh6PUHx1ZTN
c6PQcCBXy7h2+H1i50tUrEZ4I685VoZsQ4tLRibImUbY8eB0NTYvHaB51cIR6jXw
tzWxcbAikK4I0tQA9npLMLoUisxk9YwwnaSc89zHnlGCOnRcWkO8Lb1XtdYVyv/v
cySyMFUV3N1Rz1PAUW3VXAykHSSCtNc647CTBS3a/CMPmTJrDduw3YEAgBnnaFEj
+FEqf6BaPvDeqwCsfg/p2v32+W5awVQ05pQ3ZNQjj8t+FyISbWGWrCIX6B2pyhZY
lkSuO+k9lftTum03Ir2vHDrTZRR9bQGXiEugP5PiAA3h3Kn3OgOLZZdMzBda0zMf
l238YDN5bC4maUwuixL3Igmklfjg1/+Y8H4C1+cdDFU+o4aDo63n5iHdOm+oG4a+
mfJ4+YPlmh9ykNoZCPKbfg4NNBE7+MSciEp5iJLKLUCvlir2g1k2KSJlutU4Gh5y
yR08tv1TN+2lid2ygg0t8loq2jVviH2vQ3WgPjUmiyPXdQJ+gCG1k9LgPzfwZrvd
49HPp3KyHlv4qtuDChbnUROVOW8HAMCFGqhYxBqbbVPrKBERU1Kngxd3jk+iYoz8
mZuwtVLZPBd7P0kr+IFB+LPtrC4/tyNKyp2s+5m+yT5t3M6X5Ss0gaeY8qnbplmd
6A2J5zr6c81kETM1MRoMC4ipf2BBzucA2Li2VofnXssUpMbmNBZrPvMaGNuix3cn
KceUbBB3/IxTpBIaE6gmFioj2wnh3aaYmcJsIktfvNkPvnboKk6K4WJmEk9NMn88
gZatXJb/sGc1E+ziSgf7K7KkRKxO06txAOCrRizPuSC3FEem1yzlNNYmRSF+LdJR
SlAQQpRo8htPYsZPz1+Ch1NwGVVKj4ZqxaaoXOcz+wrVMnNU47JoIlJDh2tGwtYz
kDq9LdiiFRxmt0elZMBPC1i3PQhMY45lDhW4rAhl0eNW813uaEJng2JsR4eA6coX
ztOC3WYuUtQ2OLPxHtJMe+6BYREk+QN/eAIZhKEDM5R7YsII6v0u/V/PKDc6Sh4l
b3w20KUwjZa6IosF3EGMvoyYlgGdUGy3N+zRf55MxgDGr0v+tUCRlo+vBgTokWmZ
7se15GAoC0uEILWNgxbF+STPGWYwQztS3S20DOg4+SSt5yZA8L5kWbbts73Rd9OO
Lx9p6pxEvE9CR1CGAYkJH164oE7n8l0Hc+dcYfPiUiJIlv69AAh5jIo0fxishpvK
63o71FlSU8nMdG0YgLbUTY8WHryTxSHl7a+CAJGMqoTi1TvfEcHNb8HU48x7kCMI
mWAo4wpnzt6ZVr7gZ3bwqrc6nq5BQwj6tVKaS0M47M+74GCgME9TjQkgoSW+0ZaM
QcSPBLaTEQAA4NVtyXkfgi7WIgpX9WvTiK3swrYmRQIXcmODKAc0275TXLWMtTl0
MusE6tlul/ghn6+g+hUNKg/3ak4TNDs4srTHLa54WWvcbCp+eMHT8NA8yQcA345m
pMTQz4tkvnToLPux5UY+yolR/Vst1xUSg9guIpqCej2/L3eMwm/lt0xclNYoJDpJ
PfWxnikdYDbkwGWTm0g/atfLF4ptyEE7lDU6iXgSYPR3mDuxHvUeUCRMN+zvrNvw
pRNn1lozaC47MDng/C0h/v/PhXfWxcb61cvSsNgyqwrrOtGmikrovDxRCoYqQ2/j
gzfnkC4WQaUjaTl0PvTz30VD3bIg+VW1j/PXmeAQ7kHu0Z6KZSQZUqXwNZLThPRd
uMjl76FHFQ9wQxiIUqfY/90pemMOtzvo/SypNvNYfUkLstN3a99y8K6NX7cI0XDL
vC6afi0FY44cqYnfCNRIIfGh3vWAiRdxGfEpqyUK2sCvN4SZXSnJM9/QEPxEWYN2
mpWsbmYNp1RsN1CjLXcZ1/32e9lDbLQx37z0u9LlcCi1feaycDLcUN3v8+psC8v8
er933b/IA+9y9Gn1xsHY/knWqQgIUxNPUHuoMp7hzJ+XWMPUZnLtBS6AgFiCVHYa
2g3r5tYFU5JWQCqKVLiClTiC+P4RhibnzvUMLUiiBFmEfe7ggPDumJy3jZT37Kq2
iHZYyyH2mMFH4BL3maNsrZpqh78dI+JemV8CpLL/UPnAjVOULU4AYJxwMsaJ8r8h
HKcq0Nejv3OMbSJQ7SxfRaOl03/ibKz2L1tKdvgHAvImv2+ITKbjcm3WJx3U+44R
TZVs5WuY2U8y3eLHECF5isa2Zzvswe0RVtoqNlfbY3nSSXKjpziU3fWB3v7lc8qq
4HDDTA6A7rur4IprBsdHXCfbtz7gq+HKH8RII/JBaZzk+keXiw2rUc5y0FFf2c7n
jWKqA/DAyes9OZ6YO/8/4sYPJO2V4ku++7yn7h4RTjVrGjuE6GZCXgnw94lGFZim
NIal4uRWP68Hu+dqsuk8VOPM4RqPR7beK5rf2BDB//ZhK3xdbYWnj0qdmeaepHlw
Glh1nnaJ+sgYkjnn2TnxOknre5p1mSvxHYzW4xnTujZdhqxXM1FN6NTx0Zx3U4St
VmH/Ol5wa6/xCLBSay5P03PtP7iS4qbafGCNUfokKCtYJYFr+QLjibUK+eDrW/ND
rLsAifcDWUMa+V/eQ+jw7Ja9f0Eur7O68Vhb6v/DUG1YXkUb+1S72n3gCB3Nhmv6
v+aPwjjW+APs8B1RMS83yF14a7ZJefUlv7/qwH+9jTP9rvd9oiDQNne7oM4cIH42
VdwTkVozaPLc0Ciz86yOlKM1qH/8gyufcFrCH4OYA/FHIwiAEg9HB8LeUc1SE4zt
79bQuL2oe1+wW+72lW2lGvxuszlQpcwXI572HSG7DnYwYOCVgdlQ5UCHf1cv5pRr
s0P1GA7qjstWh+D5dMuYzZqALVHu9w7/w0N5eGR3eLthKVxAb4yWGHzWDg2tR5i6
BAoooJ3/tmfi7y9nFp0CSFuhpXTlC1FWm+HfY+/oczjVxix36clZpQHq5yEgyDqt
Mc8thl+p5BJfs2WZ8AbB4g8OfJ5sdrvCZZrn63QQcQIR/H5fkQnSZ0yl7hBKIHdv
EEVc91lPeKtsSZTRDy4R2lxcO9aJbuuFUKJEOg1j08qrgm7e/30ymxH6pbgnHSiD
Yz2OPPsXL8d+dqpPjvoDHmLllber8wZH1O4okT3zmX+6bd8kZPy3ezs4GUCJax9l
Oo8RaDiSDpCbky5zYBh7KoQ1UcHr3BCQAh6WlN9/HpB64vmRo7+WFLhGGO7uPHFf
RPnAqgX0PhQGHoHHe3k9OMl4NFF7ijGUQxQAn3TS9D/JezItfQAgkCYre1zX9JVY
a5RBHg21P4C86MMUoNzpOwF4tlE7BvS4K/70hGJ/WTrbnmkvvizwplGMOJolxlxn
esL7z5xkhs5BpZgff/DFe3hLcRh60MrgJ8wPNpMalECa5WMp938eDlfGhgddDuFn
xgFZzd6wrDPh4D2//c+uo4SroJ5o6DlPsc9kWWKyuCYiqqyvHwrvyl8xYpkGwAih
jGn+X7SjUmyHKco2bPR82AKK/r6BHcZcg5VtYfzIJJc48zHGCVn/Xrg8L4OqexFp
Atf7KIiFqsFmEWP2PIWKDuwkEU+crMrEIKnbX/GemzHsObANxTYZpGD7UOZhiMv7
2mwPGFHP6fh4hFARp+1ynFerHUnv+Kqq8EEmaJsJHQVe6eNys5YoEYb+mniWUHAz
n4qEWPqfZuv+GEMtid46BTrmr9X/m0F6w8goouJKOEPPmaDSoz4Nj96z2A6q259T
LOj0poBZHcsd2FFcjMlrhKURY76wF1ISv2jKfdlhwnkbS6jowdzThema4ibwdutJ
W+IGNUp+FzDHBRP3FYRDiwRZDWxKx9RNncnYCAFP2wc3TVEsBfDDJoEeXQzBKrKq
SSb+9nSbmGAY9IxOXXT32dBUJb2E+5aMLIvDN46JiujL1R9GRip54LjwE5QUCe5S
xSc0cPOygSSSjBP+/iJYXBiSZRYGORrWihjd7xL5cm0KWBoRpHjkKkl1ERC/qtwK
zuLhmxE/FCxkcKEE+1MhqxtLhKG1xbU1pJOvFiktP2wGAH3tGlHuprVI+oqngZ3H
UGHilAeaySnEZzVEzZ70DkyK8EuBA5SOdMOlxjhk+hBBiG4H6fqjcWXbdxuMb34X
PZmNVufvC33JkzFpW4DtdGqd5HApnxR4hAKdboHbRBewS7o3LEp8r53D+MJzCGCn
zVnSk/ndMo+gZ+DT8zMHsst6Wk/YEfVvPu/UQen+9W+Qmq5chTbVWoYyZVbNpYBO
SKeEzqIYd+Qn9yneckTFAdlPjS2MKWqIJOVWrjt9XXuVEMqhLjJEt9kHXX0AOP1L
IULOMS+eFwrOaUqRJTulj7xP3Yuvc0RSM4FnVbe/F+EkuqVPPcGEcxAO0CtlKOi0
kZWhPIB2Rgrc6c9cLwRjGtf27rY7XyIdWLeE3jvRyyjqahj2OAL7uTBIxGmn3i6V
KhCXKzeLVagELiVej0a0Eyjh0+sbC3E1tTJhyDZxi090YOiHamFWOglTHSUQNe7b
OnRk/WKmY1ur59RwEHarwZaVeHYxNO5VktuvnWoPGUdOG012sAFIaus1kVw7pPWz
h4+tCm43UuOG6d+LEWX1ivuGXoabn0zyGVKylr8fRMHtZ5SgolSMbdp5IZjA9V9Z
DaY6iu292E58C3udht93vOVUoftJXZZK0Q56f9hvV4jsnmCRkHsS2gasTSgojBK/
QVBhUO1ADQ3eJayI02GFVvlWvAmDYDcvWk04ITRZMJxxmnNFw2gw6jdKisnGTacs
qUcpYPoV3owRBJsomaI8m3gkjRCf9cDzgoI5Lh8MczYSEDu2bLeddIMxW3HVWy0x
oeJFMFLItOMXqTAWQcbttPgusPcg8fvxRzXckmp0eYS+75IGNX196srcuU1xlVuY
NLIKIg97srIcx4FYvXf7sCAYoXMGANegZ8Ph96F+0wgkkoNJROmRnC5LyaNd09hR
k4V6ZAYfYWpqA18T5T42R5uS8oAWtrc7qb6/HeeMrrs7AQ0m3YLQuZ7WNRDBdF8c
Y5qz3DnZtxiyYecuTMetApO7nPYWWpq1qn8X3coTcsdNTRpetVI7DkIYQ416m+UU
BnosgvqvHb0ZMsQrRlzxyLc13fCmCk+vrHyuAVCIrqEVc/+2Yf9/l2zJ19uzTJSI
6oFr3a1b26EnsVqnSkD9Jqk4GbKG4frve3XGtDr/iWeVQVbOwqQc8uMYoI788hah
4XLywwoW458mcF3dGfZdw3+Qai0kweOt64ZIt8GMpakvS1LqUvmjoGS3IRzzGRUL
P+eWfo/5UCvKp30T/LtnPGuB/091m6p6hzL4CqP2Hre4WIv8UxMMImXzfN6Tszn3
KSCnWcGd57BqmnESfB2u6G1pvW2iNdKtBXXLSfAtOpbhVhGWQ36ZXwW/oYVeFiNV
uGTIXiODhWMBs8q1d/ZCT26B0oL8ZLQzj2rymMc8K4B6/7lgMPHb4fC+IWd5skRq
pNqKG63rtg/L+FOtQlRu7DZ0zImZ9NfMYsALLppA8uHFlXc7kGWLVkIbVnnwgNuI
ZJrM9TGA/09ewMDgacOMxHdiXgj+uTbzmg4Ha3e3HWMjzxmMK9rQT5+R/9F0XHTl
jNspJ1AlDezsWA6hrB6WjgT0CDqbkGf0KI0Mnr4iQ033+dz1Jnbx60kUgijqdLbw
K2I9/RWoeTfv7UZU8I0MOhxGTL6J+8P2qiIA8/VCLLPpou1Z/v1aStzMVPpUsxmA
f1XRDW/+ZS0xp5rH04UwHGngaKm2X4fokMf/Mg8weRbb1p5HLFoZBzaSt4e5MmND
CJONObUaUTf8xFRsw7FiOJOwM4F3EHD1Rb+3uFQT+UWsK6munynxMKj8Suy3iasD
rQCPKL59LAR385waTa3qYgBdsAtkC5lhZDjdCjf7JhU8mKq9lYdP5dhAi8F0tMWR
0NZbMhmE442ws88iRFeR0JTe8ogkvuNgr4kMf8nl+OA41WIHHoXLaglhHSNvr5/k
YnG1LASJLGGJMP01YY82ONyDKai2bHbraJMg42BxG4D/ctnbdwbuxLRpsbuI9Coa
EYtAgq1fcGNSbj3n9Ul25qbZ/Sv0HQmc6sQWZjRR3PXfMlo/KVxYcBjdM6+/kCaH
MuIVh/smKGoYuKkNwMjcpDFv2Agw2OBiYdGjDpPpEc/A3Ehp3dmItWT74z0lxlR5
AiuCyKM0zaFlOYb0ZFjuVVJ7UAe9IdGqUuvOCo5uSCSpXgbmhenrt3hhW+Emtn44
+jBpP7TAY8JghixRN695DchlW9NXtM07fFDsrjHMmmENWsWWNE0w0TwJV/C6fOD1
ZpIS+ou5p8HaUYoaUEkiQsfq9KRHLIzeFg941qd6FejocJ3PZ6ukDH5NmuOjUu4I
hr0nOAQ4D3Oq1kajKRWCYo9yDbqX4txulD88XoF4/1TD0Kw9IrkTVE8ZPhXnjGFz
2HXfxV/BxBZP9mFgMZoLvJbcY4G+T3UYBMoJsdHXNFZfM7v+IeKUlpuLgP8kxcuh
jImew6Mn2dd9QN3Zcw0r+nTpoy+8VuyKWivUhtGBXDTukIKYpKrmnUq+LPWgYowg
i4oTWfIKIOPp1qvuQdPqhufaEFzuz3e3dIJznYHED0FvnggNvEOHwHRJ/GOwYBZG
lVWbtPZyclsUK/W2gbDms80wFE/QX3l/cxEhINsVFJyU6n3+XUbYSWwEYoxPs8pF
IiJMNneWvW5mUJtkZMQGDFGDl2nnExdbg5TcccTfytqJxgH+Wj4TZ9s5WS/X1a/7
JK4K0kJD0J1N49A9mZGKwzMBEgdfuYw7F2A4gj9vXOPOQg4gSXbsFe19q11Fohml
2zmymYbGiVYmN8MVUXIjR9Vkb/MZy3g2H2ROTT3HLIGATqoaoxIcva5ABGUVL01m
Re7LEus/cj+ecDSXxF9ZqSCqpYrzZZok+mJZPow0e8seBA27avaNGt57Z8ogEHC9
sV+JZvEQR/qOoCIqkxGgiKu2iidXth78i+k7ZKOBpywgIWSzJatSG+44Okv2zxFe
mRcJ/WGzJ6U0lWp0rovuHT84Vw22U6tpcSmmiL6rY4rf5dg4ifN06msBQNCYScD1
4L1g79IaQecuKoy2JavVfjkuqOV6CtsEeYQvF6uhEq1DcAdqQM7S0Ew5qQLXuV9J
Om5vuwEelu8IcRqHzkitlDdpE1uaSsAypPOKm/0GbHICnmEfZfNR/DlMtaLUsSUt
9cezw/22Vdbk2rVhYJYzAp719szA2m/O+s9HyR3iyM8C06HLAbc71F/m5+1itQN6
C6ebTPBvgrBfkFZ8BKwRqefGJ+0+cNRvmP3HybF4NGWteibs4Du7frpaSQTcLEBE
MSiz9U7h7mY3m69tnGJDyBQ5BXSv9HJI86siku8+Xa2qXbjTk8LIVxTfgUQhAkkF
WZEhchijAq28i+kOkXkK/ZOkdvwua//Z9VnT/sr+8Qb1EjdVOwW9X5Ob2jdy9MfT
aNIVDNGN5k8nEeIJ1UTP5DoAaHbZSj6edR8dq/sTslZnMkQZ2Om8C8b628yDgU0Q
rnGab2eIl5HYTtIkAKMODO3pJaG5NVHL9khxbDGZugypQrr5dpr4zGPepudQN0im
ZePhIIBeNr/8m1SzNVFRlaO+GMp6XIgbj1ttvvAJgDF4ESQS8feddK8Smjnji2nX
9fZlYhlNgRzEuW9p/7qDXh4sinvVkz04bjl3RoCOFlz8Xu8gBsIGZzSL1rqLLHRn
8EE7KXVHMjo6heyJFo7wqUkBG6ANxJXcGNFcdSST6PgqfTIpLOJiL/kOkgDGDVJ/
WzmlQoBGQY6Ov/PLpORiBRfbYy4kZSUgTHF9v05Fr8wSh1cq98T5MVz+FZN4f9VY
2WsMjy+jf6nvQHfPk84bVbtG919V9AXWrVXRXf41xlbFisK0GS/kac/sr+aGTPeT
iaAsEuBjKBA703Emu/fTY1krWXravaZpuX1KdjqRMzlwzfh5e3gcFke5JmUX/SPl
lGSRFd237rshxHdEUR8rBZWO/fouhTkF8dZKOWKmBQ0Ryh+A5UeIwbps5WenvpaC
kV18MRJKCCIQ6xn679IGJ+xLHEerBoTC/AWRc6c159pP3szD7op35CDaNx/WQuLr
p0eZdzLiHoxhrmKYMB+ZaQXWtpxBgNvavs7powOX04mdZNbTFSDlc2ivnZ8idDxZ
0KVHIKU8BPGUAaY8A7ByRfmumIbolPnij6HpfFfCgkI7unEJ33mVmmVXozLIqe6C
LvJ6KFaclZ8Ap6j7eb3NzfUkMIBA5uxvPZ1i8MXK0RpNbmfXFUpXYjl46Q07g/zD
cGZDBu2bfVh6B7I6FC7h9tgBWVKzfEGBIYk80ICmgCZh3Pk0iCc2hxx+UgpPSyxZ
FGlj+L5+7l8qEVM3Ou0uhW7yJq5nrNJg+zXd0l18/mE8feR+aTL40CkN9/ZdV3ZN
Q154NxkICh8jv5DsJcCF/ozPBBiDTlx+mMMhsNtFPSc=
`protect END_PROTECTED
