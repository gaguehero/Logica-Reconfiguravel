`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3rkX2lgchm2j5ZjcgJqWCdqP0RkAuil+N1kEMlSPHuVwerrvkduXeDdlMnj05ZGK
vxwb8/dESaDucXG4tyM4rbh8+jR7OiaMRiniHdvpwpeaqEaBiHlKraGWCubt92lv
YpticCdRnW6cb+0pEiGbu79/FM0sMuiBGfKvjpx3ZmogLOa3Bj9ik30SrQx8Pid3
Jasz6/e1z1GKpwIFwc3scAvxWxheqoCdzALjrR1qTdAiVc/1t1Axb49MS+FwuF1X
EPUE4U7WcaUJ3F60ObIbmi8jzE/b56NuXtDekL3txmMK/D/+ZxI6S4O+yTF/qLdw
BGyk22UptOq9bX4owmixQuT2TONYTORnh576u0m8x2FolJWSS6mTg1GOqn+5PFFd
F03e1xGUL2elvvCyxLiqzrD90P2/RTfg+EgnsOK5N7e1J3JSW196kxMheEg3uP6f
3y/PlpKmt9kSDcy6GjgdhqGEnSMeJKhd6Ed+X7tlUNvoxboLVn26gJuX+NhtA4kL
6oNcb8kFRR7ahPGtdVQb28t7dPQqF33xO1i8pZemUrpQ2P5eSUaClZNU0s7vkSYj
OBx8NlF7tjTd87v3/VePUJFWn5mhTgGHamUL4syf46WSRGF5sG3yWRERmMBa0HCF
m6tNlYiwjPlv06smu4qdtamh3wwQSfIn1lhmS6oJKzHMJmlU80eoNy6Z0jZWyQav
NT65SbGVilKhpdIkt1oCA22JwLjGIm+EiypkcLMyeTs=
`protect END_PROTECTED
