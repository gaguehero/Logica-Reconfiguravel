`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yoW7max+vJZoZ5iWwsljaB68EvlLF5h0+2U7fMCI6LpAJR+sjzBfz+baVf/1bEUK
gmtvn/I8XjQ6QMRZann4SMda68e62Yb8K98787I07jQ2lHZ7ZWHSPYmUI5XEvQ96
2eyBcf/+YWKvYlKPGF05dCamZN2HlS+gswZiZAOsAPGkcmpnZIfpVoBCmV//EK2/
JkTv+wY0dmHyTF/0it7humb6s1h07JUM3YM/PT2MS2VnauV2SNax6MtDwUT8D6pb
QWRddFgr/7mNzb4vNBzntvGM0g60yfOGDAk0UQVdYqgVdtLBBEUzY8MYojQgC/Xw
Jy5DzybT9BwghuRRecVt1icpXw0sNm6Vf+6rUelF7tUiH+SKESb9UKmdu94gXGrx
vjYNeeVMDdIu5tJyeUJgWsQp+MyGZmsQjN6n4+Y95fMLpuPS1Rfrzb2b2e2tdIhs
w8VdGBUiQ/wAAou5QJCzt4Dj7FtHsiybdtAduuREFXQNsXmvH0Tktzbyy896A85R
eN2dT7pbpK58yC2H9Bao6FyErmtjYZ7idsPhS8Ca2c9Gf9KHfjOljnQzMLt5mqs7
5FjrsUKa57hnoCRTvFkZOAwBBUbMm0AJLYRO9Y11e3biVwu3hWAdJVbS3KR2+eM0
az3VDKWfHVH/RBeblpZRM6M6DdhQCoSeilrJFHkCi7P1yS+PduKj+pUplOBLJpI9
H6uzbQMM9QEokulKoJYArxZjLrbh6KXPArhYR3xrk/M=
`protect END_PROTECTED
