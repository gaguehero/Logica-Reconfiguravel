`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xx5oQC7CEUIH3/IVJfz0osNZKG2Jj9xNbIRHZkbz5sjrcJ3mlP7zAF/z3ng2HrJt
INAzz3YO5VpGPdxbHGB3pvmFdS+nQ/Byw/nmIPcKLKGxgTuAGHVBLXNBlN3oX3c2
m96tfcDbmVxDvudirujGK6H0l9sz6Y65Lz/XCmYUeDBduWBP6+wvw+ZDXtapQYE0
wijvzEGHDsyZ5ugue2RxGG6Wo0xn+lLnk96jcyRnEdlGKKDp1IUJ6tSf2FLq5DIM
U7rYloE6NIyofkKSPML1dKgTODHKHYj+lkPG3U92V/wByzg/6FtGWNndR5kB+DIT
9NwnGBfAKENCBnxYectQMGofwX5ENSaEAIoMxKO8J/QnEb0ITfpB9D833QPtAJjM
bLr73eAHYmqWPQnaar0R9ezLOFKhhgTyfk7qAJjDj84Fz2Icnr5/8BSDMz2AnJdg
fjK1vAMx355DjBDohWKk88ZneMq62CUgvh9GzNTK+WGVICvQ3HpWNG+lkKUlDUar
Jy1hwSgjoVyOWP5JFHiIrY+7mlUXS5pShosW7JR1SdAuORDsdk7KYt6SJwr2SoMZ
0rBy7EDGB+EjLEvoxcIpdNQcLX/FGDn4eTew/PXAdhbbvmbKhh4d2CR4iI9Gg2l6
eNmtyuc12yPXKDPVsi+UfHeovlSeJj4WrIUvJmOqMOkU2TZ7oFf8IbuXiFzjlpDJ
PLV21ZtCdFIfPPIT+Rv2oEf4Z4pL3cUf++zwoiUleEJW2HvAxdbo7poOGzlPkkAr
QHcWpcDEmP1/zmihjtkIVYWk84ICqPna2K7lj+InsGe7EKmKqFdvAw9fYHq0ZcFg
OoM1XNcirYCB6gtGheQWNNKKESKggnGDMq5/XAK5jl2Ff/DSXkUlDW8UWBU+gny2
Mz/7QOgbZ7uVcluaVE2h0ji/gq3JdUT6kcOqvb1k0zTcvXBk75ZD9Xzdm8xEJxk/
FM5xcMlwEZHQ9WVJJCe8sqlrrn3mPGFs4SI3xHgBsX7CpClbPJ0bxBkni6ZkIL/T
fFceF9kzx+a6K5sdzpAUQpO+DXuoNUEQVijQbgcBRF2poMtq1cYzG8OSk4/ORWQQ
Pnc4ATYvpb8xfcE+PX5U3GXpZf8EwQTlDd/VKJ20maARo8oOQbzjHD14IdjXmQ87
YW+Q0T0dGirBsmMx+gKxCpWBIx6mu5/8bBSpneVAAYbMbBWGSHJRTJmBUb/eM+Li
6IXj+h09t5qMzLNij2BGr7B6GxDi8Poq7YiE5KzSpxJngmnfogx3H/Oxq9O1x8kC
7+jEGkGtVM7VjJQzOD+oHDPSl4LJEaHfyaXS8nWbypFcoDjTqYHTfKec2kQ39dcn
peWLp7wMWZtSYSH5DVa0Fi2EDiXNsYt3WXvwZPWVUwlU523Y2XzW8BqICJAkMBnn
AY4IddAMUuCYvPoR/dJfrjykFphTB8ySsBBNbO5toCWEH57FiCiPJlPrRdhdtLo7
zZWv1M4ZHXqh1lvuy0VkXf3OSumyaoTuzMPNJOX+ZiHEELuXYvtZyS42668W+nJl
1de7Y1ERnYcVzSdQX+EbaCrpiA8q+v7alVLPX/LqOOVlwBn2Cp4Mg/MkLJZZ2BZ9
5or4ZO9An6wo3YobkiPlrW1XU0L6oVzVkMnBqplDHdB+pPp1chW71N5eT24H8az6
4CugQDPIS9SGw/K1gDasOzFfsjgVLQ75VNeMu1ii2SXrpej+ZeVaBvr/ynXYowC1
ej2ENdNsjMYIHrEWTBn63L/Axe63jXsgaDAv95DJDhG1CjrEZ6KPGSeIctNNXrvQ
QfBxyA5eckcbHddzEMhB/cyQ5hzmxSYcKB0guLKaMuLUkpA4kBj0TWgKp1/HgQ6W
ltmTuQBolS+kiNpqES/w8n2fXXrKf+6PR9IPoa5Q+Lv9IVQ2w+NLZZrmeplL/PAG
NRdQYT4RT/mlKBWMSNMcs7wNc992xyE0Qie2719/PWTfAEv/JSSdwJVcnLt7NTH+
x9o/Atssd5wOiOAatgab4XZoMqqqOyauYe0qy+/c6byexDvvMicuU7Or1eO3qdBq
cQRSSK3wrYAboGRKjD+ZWQ==
`protect END_PROTECTED
