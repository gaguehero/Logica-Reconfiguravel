library verilog;
use verilog.vl_types.all;
entity cont3_vlg_vec_tst is
end cont3_vlg_vec_tst;
