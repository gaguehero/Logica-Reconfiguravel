`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGA3kKV4uQ6NuT1YnsJxDGc/o6UpVV3C3iHR/+0yuQMZh5WI8kazktDcOnpbGoaL
KdCXZNAt+mVV8Ezs9/qqdBNsDyTYNqw+BbL3pt/JBl94D2YuAZ2BCCK3jMPXQH/z
TjopS3H69tdgckiVp6h55zVCEpP+0ST5MnVhQp5kUs3I4jEMKjaQv8FyoOVjRpot
L7wREtWZeBdMRvCsXekKbzVoepqCepqxFBv+xSPHPLkgd0SiW3juf2mSaaUSz476
E7qIGesN6na66kz22VpiP/EogGoG1ed6TB4+mM9xeoX29hZLaWL98pC/XMk/+Hme
ZNLJf68ytoiRtA+HKHcPsgqtUhje/leivqMuI1bIUlm8+oxXoQ9ts4bJy/kr1oFh
lYPV8NUmoEs1dg/ugcz3H/5Hx3FqnkAlHWgPYtuD/ww4ANS/2rqdOwOBpc7okNKu
RxKB62FR5herAc9/bMaD3wYmMBDHSIx5NPZm1YGVSnp85Rq/CaJJOuGugM9A0QhW
5I5jDA6e8DXwLauixa4KLTkz0LbH17MyX+GmLIVEOSFGnwMtbKmRxTNs97/qgEfw
KKf0qQyOMOckyK+D/7fsrwKRT3nGoqK8fLuOF4CWOFoebijCpZz3wHNVahm1IV1C
P53tu9XgwCd62Z75t8q07uDdnvhTqiVI9lMuEkqXvVflcSlRyprw+zX+Rw4g0ljK
ewvTYAzBrlE1VmmaRlY3QwRc8WfmY7uRncxk8B0WFFlc2ymrTrAEICT+afvHUn56
aRYAO5ZmeJpHxv1l8DsCffVIOJjJulZGMt10fqX3MDzA4Q/BXwg9/UJPsePXrM8s
Ves4hGtoF1ty+OFJwAT47hSzTGIsrqU5AxD97QG/1DU6NWvNpmue8QE7A81ftlVf
AKbd5FYNcaT4/M7L3Fgamry67CzP4lmX+kQmT9F0k9uhAE5+xWqo/bTfNKax0WGm
WNHTPK5QIdIhuBt/Ex0IVHOBaVmC81dh7HL7B4Y9Iju0dAElelKV07OOiOEziBs3
fnx8cy0h3XS64yqSjNYozGqBxwqllfRNKrGvNdk2ugdb0LxGMs0zmvUoZrwCZxYQ
K3ayrHTb9nEV/OlKrO7UvvQABkOq1ev4sauOqFovHim/886DSi/7csMU6Xvrso4v
Kv596E5mCTIpMSfDO+jvJTUXZzmT0YGTHE0HV0DDmdIqVMtHnj7YuaFCf3crS/Bc
y0kooF5a8Wdng9Sdq2pIBLI4pp17a8FmkwY21U/69q0ItiaZlBS04RmEO4QdZ/yt
Bp4NDaHQuyPArP0IJ4GCsw6xUGdgdAZtmEeK46qsRPLl+1L4Wc1YkZlO/HTzVEUo
CcYP5gyGr2CFQBz7cY5dRF35PYyFo8zTUAosR4rknLyTXErIh/dhfNNSxRTTOqq5
L6GPOio1xmJUNcKzwQAc9Q/A2bDiRcuMe05ZFH4XY/kG4xf3H9nwmns/s8ZUjpQT
Mw9cCtmjCAKIugWt2qti6LlMGen2z9DZ+GyJlGbA1XWWV7Gf4z6Xzwq6Tb0K0MHC
vl1pXEB6J+iWe1HYd1UZoNrZzP7FSaaA3onFxCC0VyHDEq1STsRDAASnq19Xyv+Y
i2hIH/11XQ0J2XKW3t4Xn96X3faeMa9sLVZLgeg5tSjTUQpHB2+4KLu/s62bCR+r
4Q7uaIpN5fZdHxAxk2kGAVvjiY5wTmlNAQfPC/dRhHFGehRLQJ8Rl90MPcydths3
HgRtbgKQnN4uS7s055q2zSgqkUqwh+yYkaB2QGD1dXtI4W3SDknFlXpJwhgknIUM
dEE81QWt1JPVnmmbfnKx4hFZiSYZzunLpaDiweu0CxYvOGlScaUH8pdVlG9ZbTvg
ShX7eEWKY46gH7JKeI3iEiOZIhUruFQVwlsjoSWcmXKld+OlN+sY0PBuJBOVYGvI
00OK7vCgaJKNcpD/vnYSjQUAhqHB2pBfNcc8Y8nBp/dwbfxyit7kqS1Y2jSFKJBU
2EEd6CWAFs+oUwfwq8fnx1Wmuj0jc9avTzD0M3Q37ljr8J/Lx9Vh3nNc005TY9Zk
`protect END_PROTECTED
