`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6AopNrSnTro+/tnuOiwEhDw//8LZL+V72LTiv+sL1EeLjw4oT7hdVNZbOgTzc9j+
pDXbgaNMYUNpmMlgC5bUUVlp+5gVGyBtVOvACk1A9hNzQWNPfNI8b3UknRzYPCCk
2xIc4rOyDZHZQCh99eb2kRR9MzSIcxg4W5rfcEi3gxGFP2o4ZSQ6zeFuM4Lr9Ogt
Rx7gmGn6RlaycES1bp7hKxnTPg0VaMkBVWSCUNNmYON4i8yY+J+Cmk3BQSWpemE2
KQ9K9YdiNWtTkdzM46adA2GA+aRaKUuxhM0efhp0Oo/+P2uPwfFzNVOz1WzqSgZp
9fxw9UANX28uYSos/fW8hfS8M0pyjFUFEBNpMH44xp1EWK3ubJwD012bmZv5x52K
VYaRa1r+oLv5hbShd+pxV7fbV4Yhch22d7rDlsRhEZRdEeFfcI7HOlWbLBxjJdaI
+lxwY2xmT+C8+DqBplnc0tnK2w3Iqk4n8MRj0vrTCrekvUx0c4XVbkGiJVBeEEZs
FhTDvoLeZ1DwJmZlIaOZxgVtmJwH9kR0UJeOCnGUBIXFIi8SASUXP0DSBlHN0rNf
tBRjLGVUuf/+9LbahVcRE0KrNNJNReUrmStNL1M7H7LDmpPHE2Ouikgzz5RW4lkY
ftXZ4SRr0f+lx25i4RKVA0azcOQzyRf6QtqfSHHVFhRyj79B+sOsgfvi7o47T1n3
`protect END_PROTECTED
