`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEBZxnS2R/1pdjNgDqHJZvSdQlnECD+KvcBffkmfFMMo/RPLHwGI1+cuPhtF6QqI
R/hXQhLkP1I32QYsctvBiqoaJUIeViNtRBRP7fL6U8aRY7KCrzqNhGvQWvVohymi
Q0SUPbMZdwFfBNyQb2orVTGGd3OSwWq2oNOAJJiwKYJQYnTjRsHffXsKxsVdl3s3
d6oGvNPSY1VhbfX6vpDQ0ItdbJZxGI2HE986EHk9VXpy6JAcEDVX40kJz4fa01c9
rOQ3u9OuAuLpiqZrL2zwa4X/FkQoKRXUEVpSFkR9pPttX3KlW6ffTvch9wxqnzDH
/RjpTzcCqgfig33Uro+gLnkMG5yRR/DzqJTpyDcs/sjYwJP1P2jVMXrcRpcFpw6y
JTZQ50GHuoeP5UCCBVtxc/HYCLlSXpipOFRHz70UHH/7NhKLKhG2s1u365M/wQyG
K5NdJvWsAZtgqPYTBVcwaxwilUXtiZLQ2yzfT89pizSmE2J5T7xKeGRELfT92V36
wFuLLT7o90/mTYPa86CHc5rlRYsY3bJcGTOs5tX2hg0yvRijrkLLJYl+vmpRUxCy
Gsq02La4selGG4r51QkUxYLJlg1d5v9XfwJmKhgmZcc=
`protect END_PROTECTED
