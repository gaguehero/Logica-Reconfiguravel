library verilog;
use verilog.vl_types.all;
entity unidadeLogicaArt_vlg_vec_tst is
end unidadeLogicaArt_vlg_vec_tst;
