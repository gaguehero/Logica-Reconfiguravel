`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glN+xmwyEv1uZruJiTKX9t4rm4zK2YJauV9v8I8SLHF0rJTaxC3XbaZBqIRH5zTk
OxXlhtosIpD2yV1mjDibtaihx3sngQ6WCIrVZqqTFJU4PlLdmweK51TH+7fyrhJc
EvLMFZMOxqQQ4NW9qwBE2ZhjwVsNDI1vfx4jOGxXHqeGB+T5ZJ416UdCRtjKns0i
hwac4BZpKzOc6/Suv66p2IiicThWyf1KH8yyXjMJ4lajbc+/08IypHdI7uYeuHC3
Pho9xlo59BnCERAu6u4mAfpYvZ6u6+0asCLBBmcmxLHlVgL2tuqeSYx2edOSmej8
+gW/3y8ehjsu/N8ByOSF9EhpVxXKchum7iwk+7r9g6GJE9UrR5wyrMyOyfG+QZN5
7/SEXAaYz0SeCZPE5YZb55g5ubFAtYNrOZ4p2UqEZy3QPGrXfAShisdc5O/dDFjI
WoSoESK2mauj3WlpbOJb4MKCxU1bqbEH/jP334KgsA1SmtKLeM0/DuW7aXo/sQpE
vXwoZBEykwCG/xqSxQHQCBNwdmcl6rRfwnGoA2OCCiShBpsxUZDoxlkHGumjPrRu
KNCb/n4mmYxDxjTx5d/z7ZiaVqE5M2vDjH3wBAcyNLZyufhPtUQKrzipAnBzIX/4
dDwmdcZ1FEcY9VzcfbGM0xF82fGpuWx4K7siVmr1iKiflUKM9s2IPn0W+VAiJWDo
zfp1/uS/FU70cPDhxq66PiYpV9fxiwojHzsxkhOXkXu1pzLVTK4f2rW/qDLin/Bl
Mlx7RoWkT3VMVPxF43Oc6uqXjchWY7UGIbiTJJ0BukTh2C2jvXQOLst++IVzXm59
WhsVC2d5vbRcic1U0htsMw1SyfhoulpfG1zX6Abmg0H9eP5C67bMcuuvJGx9QWV0
WExLPJMBApa2AAbs4DWw0ZHyNzzxR0uf/ceyVdOpAsy2gA3/arz/iyGIPeTBuLqF
Qz6n+gPha6MjrlryHIg6lBvSFeQ4CNRw/Z17zSLdRm79AJPYJmn3HJDRHCHcfjlG
OFPNNU9M7+DCs9WcepNieu/xGTSdHi7XG+HGWxPry2c2xTTPTBhhP2xgt332uJ8a
8k+R87lQolr4iP/btIFGMpYbD7h7MwntH+5MluwdnHGXGyvq/Do4tt1QjAd6+enB
pLsMHz+9FvQm+lQpy6ezuaonUuemhste2eRZRR4KY1OQNOXSt6mFFXB9ekN5ymyY
7AmEWc2t9SZ78YhSha1eY+ZX+/j7kQNGC+Rc0BxgCcN28PCXl3FNFfLezOyJbxnu
LlCilwIfvpL3Reh2KMl2DhIJbMERhVjOctLPZUD7+0uIo1kGQ7unr/PT9BJIhiJQ
hqMoi/dEPW/u2DSWXNFR7vCX4O9eKTf0s4LGm1W2aBzpKqGAlNF6Upwai8Elnmf0
U+OHrlU8tTF24bzFaD1XPez8QXVZZ3PnN3PyuwDGpJeMh8LpwC88knZ1eOpGDjvz
nKOWEKcwB6gWjSSPxoxlOVJKEUSql226OqiCyL/fVj4xYoYO+sVFnJ9B1XIsv8YT
vmcVQQW06Z72eQ8ccpMJ9bB6nCxcoTVgVzE7oyQuSf0um51XzBfLKVD4qsLXrEe1
ANjIFhs9aJt1vv9vP0xupkYgmd/Ip+H0Zx7N3TqamXpfCio6BPgdrlS3Un4RnoPV
EAdso4s7dwP34MwoZu0fE9Hm2aNOQMPqwng6a2yRpBviBhmgr2lb/1lIku5xgNC/
5da7TYA0tnSyy7kJ4O3fN/9vYHlREG8jV5jHjviRM7thjFdLdErzgZiRvacCpMhM
cRh8cvW5VApNtIZwQ+zby6bQG45peAyw0YhBify7wGDi7UCxeEINxzk/HjnY9qJM
yUF+YiesHXXBcgKq6k6B9rzqfGbSEdHjm1Hs0PybtwQbyQK+w2U+5VWCXzzkcwQD
lg7dGYdZk6PqwjoeY0qLnEVBZCZzKw0SQJ3QIqA3N+pIArBzrllAAro+EmGTJtc1
8AFoxUQyPIlsDOMzucGdwjf2cobhFWUvM9Qf4f6yJP/TRKHc0CogbYvtyjGvM0Ks
DKITcgMbMZdtfCdxHhrnjrngpXsgBSkkim2XbEYPqgcLFiZJzhwPcLcbq1I2vBYS
1OirIEB3dGINp8xV9pP5u2qCyh8EX79fAQzxncgVEjpHO6ZdSNBdfff37TxdAkc8
Z0PaSBomOUjyYEBHZwLTbwYIa9gXwRAiJc89zoccFID4SPZP+9/qDQPC44cmTJHw
j1YhA/WK7yYn1ARGs/Zdog==
`protect END_PROTECTED
