`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
de7AY8yyF+FCNl3D5HrUcaCxMoBcr9At7aYLnRAyhMw+myNI+z4bhoaNxxKxXwwu
ZjR6w27P0OaPttIq8BF525gpCTA3BfYjp/hSRjNrmA1SGZkXiyWOWECWnpBrDgYf
8Vd+qN2M8OrV2EbFphteISgMK4EC5vpcaibmxZnk1Sd3qZZ4h1p2GpwQj0q7JspG
C7K1bm4iqhsndCJLO6G9Bd7qTMRwr1UP+TKpb12wcHESnLpE0kiF0odxdLCgFAgE
4Iw2cl3oo0tZDJjCoMkWlQJtD1Spi6GhAUXLj3z8JbiErZPa2iKTxkKiFqeyPJCA
wqVSt4hckzzhAHBFCnTSb176ZPIy/m7VgVr2+qg2xhqp1yOybqg79VedWaWeylq2
t0atxjddx2g5vd+TvbyQbqft55Lh0WSn65h28UBZZH30ffnpk5DucMt9RGfn0EV8
vz7gKbTXU/sqs3hS88BGylfjtndOQ97jqBUYuv9JZbFRV+vI4F431nmuQm3FXHz1
rB0wllFRmquPlyMyWq4xdq+xFNfLdkoolcfzGtTpaQIIi+14L5Zbrf8e5AzfESMp
AS/iJ8b4tFtY4IWasVNUhnC1wLOeZ8f60PTAo+JM1Zk=
`protect END_PROTECTED
