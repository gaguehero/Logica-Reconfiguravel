`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6swNo31mxPj0s98QNOAxHqq5TqYj/HKJO5ZcjSHXth31riscePoYbahTVPYcy02T
6P0TTM/ohWGtXxIZHTWG+qZ5ijVkpMatHLNWwFZ+cgbY6A4KXlPRZrKSp0ZR7oHP
XexrDglva65+/Aq1mZRrcg02HQK4SGbL0xDkZiShsWhib77OFwsndHvfreGfc4qt
0zneeKJHmPwCcJRh1PLUOlpzKd6kddPbtKq5LxaoZEc7H9I8OBliDudr5oOot/df
2RTPd4zQaU67sUhQFObUMjcyDjMdJhx/FP9DRiWfmldM+N2rHdaUPQbBbXv3h86P
Tq6K4HAsoR3Y1uYnbaWBjxkk+gJYWbm+jxtMNBmnYoDDaBn3rqJLrxLE8enajNg1
IsWbJLrAZpnp95HgEtnbyCY9RJmEeFLPs8Ncphh+shThaf3iTdrkP2UJgjWdAb1+
85txXWk21SJlYPLXgIy5/rXXpOfZrrgd0sUwNxfNgDWOdUw1H4wBwWUzQnu31p43
WC3b0uFwStWQ35bwhLZnJz1wIG9Q3xjeTWkLYMzR9VFVg5pquLCWvntVpYfIBKMe
ZK11N+SU7moU26Pwv8BktvuCPxYE3WAgfvmKTeS1A7BqZnjlweTHMKGlKK02mZw4
rRdA/o1DidYTM6l3NLlMWwcZCsXh6kStLle/8MNz/yhxDb3X+BiIqwqHjA2D8rbG
0ImczvGvZGjmJKVkZferJDoImbg9+tEnvCelP63jJeShY+Et+5X9NFLc572MqVS/
PbwQh049+4YsuLhFwAOOlnXOBmhJdu0ESPmGEjoLLmbG0FQcvhg5V8Uhmn6i7F+f
1/3ErgR2tZlyISDaJjCVH7fbsJQnxWidAnLQAyg5vxZKWICZAS89QMfD/IqsBaWT
rR/udYMTne5JnkmxcUgB90LNIk59rO1xkcm4RYv3aGyWvWNaHMXOp90kTCbi6GkQ
DJAWe9SGgN2C37Ev2Mx4NmiqjyHlEhYrDb303u+jruW5n+5jkdHquS01vnMvH0K3
wFoO/Ap9KN8kHQpU5tQcOddaJXydUWzBdDNGn2kI9NhHkHMLrIgXXThg6ZgzqIr3
cNeCS+8s+Kjkxa4dtSOeBcDlMKpoIjL60qS25Fe1zWpp6j9iwYwX7aOegPiJS/mF
Y009Bi3e6iTjd6+kcridrJuJkMm3X6T8bXbcAtC5WWxEdiDSxW/nF2+JJSMSgBZv
3/1Ygn7UpcrCfVY2ld0lSU6iPiZKGCU30KRZaJvgCRqzYjZUtNLQKsOGNgZkjEui
P/h5R2eI/vC60bUbUipSONihSiL6Hd5pxYGY71PFEtq1FW27Mwpiye64KeXmJtfX
y6i/It/9lS6co3oWxZuKNwV4XM/k0l4jZZqTiBKXwbcV7bpFYKB4v7Cbjz+wZECT
2yGEJRNGtFFQSTaO+IqcobhHOz4P02kUISF/HdNdY38qJfIgrOVTCNxmZO5Bdoqg
WDRMQWm29quy/ulIJDX2EOFdG85pu65NNQLX33eQEnmtDac9+GbMT8prcj8HELMd
RLntSw5XC5rOmqTbhSOi0fIfKDFyLtvTLKogAcXNZi0jAJFvC/G9lT8OrvEe4h3X
vcmB3uz89MwDqwLvz4EErYWyLhq7h09oPhG7yqbYlXKAVD9FbfZTNCeJq6I0uBwY
bfjgUvc+DG3G0thkJ9vhcHF7FJmDiYKypW5IqMpFkEJA0YG6bonwGLT3cbHKzWKg
EuBZSVIFYbuRc6En9pXSesTzDBoM5dlorbD4fMTlkmeJENJe2JmjHQmkMz3ZgGd1
LBTLKEuFDjwTVwmQxRAGEh5M2YriwiRri4g6n7EaUW3FEzjDOor8QnstynsnwYNW
8rxaiGmf9AGNRdpqOoMbYz9dFMP481aw1P3hOaFYeJwkXe1ifqIJGiGUex7TcCDc
X4olmD5CWoKszpo4pUIwpxN78I/NsgJVkIaT/zcpGusUDtHmY6OrazUbmj+q0sRC
pQ4l5Y9tkjRisJiJOVqTP6TX8YmrOHq6D8MELnn56JFnsF23FqSg8zkJ58dMfenj
3IvSTygxDy/8hZux5phIaKgptUogwqLVbiS3PTbsGIozEImn1uw/qeOTpDYwv9xo
S233cLU+eRaC/wTCSBNKoTLGszNqnbpRzi4znYfL0XawBpBo+bYdet7t0jO7sEIl
wCLDDDRBS8HVtzPBVjZnu0104JdZh7t88jY4WF6IzEh22SCmODwnHtNnKFpmXOhy
vTMjekyk9+BVAjirzC+jYP/hWbnHAB6O2s+1GPeqLiuv0YIfoUHi4VtgaXjyOudn
PWv1063QZV0YdPaNe+XlNPCCFwFkVwaGaay4FO+AVCGZ9amyO9h3j5suZo8wczK4
ybevPGI0uR5yDfPpJNY7uEfKcnh7XQPMPWjWJQizp6nx7iesqgZI9s68dmX++g0n
RsO5iOKyHIrgSeAQUKCUZe+fem+g26yChGPBaQXoozW697V+0RyYItbwVHUsh+Cc
gRXmMxLhLQOp735FhgK3VhHNm7X+g/39XPKyYWlwBwu1WUPcoXy7YP3U7uEDQ/9A
vn0/7SZzisTU+K/VvWO0Cka76SpXVMWOH9py36atx0u0A2ofhKvmu3RP/eloj+5Q
SbIdF9cU/GvnCG8mq2MV/mGjpSaEVfC3EJAqmvdA5UzOdpzgKwzxzTyY8RiCRQY4
Q7CXOxZNe8ZXHzC7U3Ij/99y0AfiKU/9ye9an9wH6M98gG01Rk9PjHtXomGZFoAT
oegRJLzCpxN+jgjr1c8l87Ff57KD2MV4OiyOyCyEOzRcV/Tq++TKYVFm2PMKsHim
Mr/KqHpPrIbwezz6QtaR8Cx0qB4HSjbRJioeviobShoPoayydeyw/KIwslhRogpc
ebhhyS70NtuF7PmBVEAvhEGrU7abu6V/Hnk2gemXa/2iCXhDL5WCiKFFe8n0Kac4
QtpBmMtLPowoKx7e89R9HTuxtj3boAmdBX3JzKNe1fc/qYtylAiu0BWjYnU8Wn5Q
WiHwCqCyHMr3e4ztblLlbgCxAKdjO2zTmonaJQ+/2lkjUIGIiJnSOfe0aDocLQ8l
PU8LYQXtQgvDdOp9aQ9uH/n/uFYYUIX1UL/x4N9gQcEQe/yqxsJM8PsxFvAUNkZJ
7hm0ltYMsOsBchZVG2Q981ncfkRcYjRgI4YiWnW4Athb5I/EgS7ODM9sx81G+7mv
zpismzjf6M6HKEnvUTijm7p8IAmKY285HCysU/wAdHwHywa5XVSr/2KpIfM4C9Y6
KaPkTfKkwISdqTu0XxfeEtIzVLGykQ71V8NYoKz/ndmLulsV1c3oJqlCM6p60H62
Fe787Qb5C4B4XW5jaO91mO/102IDxzKbvSssGQkZU5+u8kIF/UoSS7V/Oz6wYjxY
rofdhIPfGZn4viB0woJWLMLloE3ookL/3PB7kwJoMeCYVaYGRq3o5M/aTvvrylrV
OcXpSoHQgeBQ5fBblAcaOcEC3nulmMa25/yM3IX/KGPlCRNo/lsmS/g+3GaUxWwt
XlU6ZoeuUZXfnbMC4hXKPsNTWLs3/o0sXMKk4j6f2PRyCduuySqqUOPDWQX35izr
ULDUCrKIQYfHn6u2zSsdWqbaUKQaTcXRPf+MPHU4NRDXoxk+2h4iXAMQQaBPB5Dy
0L8gszogZnjHYQr6nsyw99oKZU1j/AVut/DUJH/bt3DOeCmSNr5Y3NjWxnBiV9CE
uYJ6g175RMAHRd7pssG/zxNXaa8IGRg1t+TNiJOKttAWj1iOig3CuJytnPUq5zGt
XPuTTKI4xYAXe21bzcsw7ZKVedW+ojXnaeivksgsVVy+tBx3MKdb8Zg/G0Tp2eeJ
512LTgMBSESpW2ISzPCniV+JiA/olW2Cw6ppRN4hQsX5K2g6FEDkg7A7PgSHfS5d
26FrqBp3ykdL5HgkMeDYGemaqvQuKX6P8brmGVoQKnOr5/iMTgqnMOb9SapH9cDe
9qqNFGubLsSza/Z7q2umgURPN1UbjYq1Bu713vDpzLhmoLK+nBYYC3mewJJY6rzG
nr1AhDOWAa0BSEx9sPQS+75F254Gxgg50afvw4VwwiPvOH/VNaX7WMqJeB9FSfGe
Jb035Hvab+JD0Hgrlsv4zL2lx3daJPccF3Rj6Rd8SdLhzTPg/Yeo/7lXYUwijZd1
XWyk31OukLme08JxH3pJFwjf+Cuc6CwOhmmWUAxIj9s+YTqPQp7XGmxx+a+VD3jc
CjbLtakpv1Xs1dfKVjOdCamJbRkjk4zbn6Z2nITG0VVfdbrrAYE5yPcfSk8bcxQO
KbKnFNBBXrc8MX54Puze6Y5p+1Nzz6mH1GUdbKCc1fKNLnJQZO4ILh/QdieNxagh
O9Uq+ndh7NNPWfSH6fF9FuBCsJWEVoRl6L6wFDNKE6Dq3By6GuN+MJD6WXSduZCY
hdLSo9wZnAKTW8vw53dJCp/MAdh5pkfmB8d0Y63Aw/vQeEHVipZKoCJtVmHiLMgf
v43d8s4dKqloBzJQgsSVATtGbgg/fyCfDneKro/eeasIuM8RQnz+gsInRWXRmnwy
uhcnAi5ndMfuMvUkziIjNPvgg6pHR6gWGagtGXUt47GLW1urm/eorKnFkwH3k/Pk
n7JLHuaM+HaTvmdqdp0Moca+rEKfngjI7n2MWTF/NrZZes+Qt4a44g5L6HfyJlv+
p9wUJNvYiUa0ZURdWQ2BmLHWe85hNEi/Ib9CU9nVEYNOAUnxbBo/D4jFRfp4QcWY
NhhVusLuovoy4miWOo9Thrq8olBje/8px7Xx1SwERAoCp+VgGLTJ2dUElOQjUFDy
jwiFUGimziiizkxmQPEXwxXrM59OqiZO+IDE6QOXJzNdQUGHJuNvKdq2s0luIQyl
D5JaO4b6XX2J/GoMKFN80rhwoMId/0hAl7jqQbceBCQjaTvsbBKW1K27nxvK/QSR
3u+HwYCuOE68HXTO/Oleopcsx5XHjodEVJHibitBgt7scRaSPTFpONy6inGuCP5b
ejbh1k/MHr9XvegzpxE2Kwn7e0IR7T1roMEEUe9eQjO7L8E2Bg54k1bahBnySiWr
bhBZhHwZCMgcoKp9aY7iqN3YxzSYDUH0+u5VdJ0wXSvbn+PJSxKC5DAtCpe/Fg+H
QbE8X29JGrpz1LxCpSVpDm2Ip74MNPjiJLjmhloDl61oCAJ7ROb4hswuHIYEFCqk
dCTyO5rssGmo5a/UaRGNbXj5Lt+VnhsBcQp1aG9lm+MXJPthyYWQakZoBoC50jn8
3KPbupC06a8B4suiexum8YQxzQ3kdDU4fzwk/BqNwkEDlEkOq2xuMxYCasmWr5Ly
l+ciOj7phzY3nNoL73RPWDClvwdLQraxGtNjNkSIMk4gocBoNjggmkkGIZ4/qLHL
zRRH2UkRgvPKIZE+nnD/Q9BGZEM5BHqPeNGjXbXOpkpWCu/DpdcYZpwAXF74w11m
pIjFMay5HdYRsQUKKtdw7nT52ABQep+g1CA2GQ0ZRtI1hbhpEiw5z9qfgiutUd+o
Tt7+ehBYMRoLUNeB7LJF6l8rUDzT6dapBU4vbvICQAuVLgbEkQ0KydI+z4ME1k89
jyHkA54PPp4MowTBoGElZ38P2GYAt10c0B4C3sXdek9f2iMWvloaQ3JvcQ5nsXC4
rkme6/2Wygl/unvvJ1w/B38KscM253GB1rgdjCz8OPtObqtM5gSVagFCYL3dpGBe
cDXgIkjqSJXLg9mho0m2DLVDs+2gX614Iaf/OEsdICaBZygOtoJYg5qr3JOv389I
5aJtgE1VowqRqYg25CotWXaRkh1cyy9pasp8CPYT4QAnJO2m8lkJIfsBAdc6R5AR
by0UHqiZuYkKWE7OfmED78JPMRgN2TnhgrSFsxkvuNR59Zsn1IoRIfw+Mbvz56XM
THLV+Wz+3Wb0pwbBGkGBdZ61GOhorcGBArk9+TZWDv6AoyWP2wcxx9ZpDilKBwAZ
CfvrygQQ40cE0Ygd28jKCtYl/UGk6v374hmejerMx/lSGGwBc4XYurhBKMfXANJH
eOu0C8JMy66DLDDDNb/VcBI1T8yFAPHpvGQWVGuDIQ88QVK02FLxxSNh9VrSFf9r
MF2kBEBCJJm2gRrvWuhS4b89xGhqX4MQlwK4otC1nm6CQ3ULJgHIbHdS4xLWrnzi
UyxPmWXJPC86fnYVM3nkekfl2xqWee7BmLpSK0dJIEvINDRQIYO5/ZAB/j+ch7UW
9WaJhXz3tWcnrRwCjEbDPKsNLSETxWTgk8WHZ02p5Ea2uHk9uP+jFK18yoMgQCXy
2IWAHPJWnqvFcDbSstUnGmTv5zi09i20LYFRT+HS4rH4wqzawkR5WWjRF8Ahb/nE
liqRxERJkg+JDQyTDs6/vwGDjYhiOIwygnqdZNo7m1tOClOqHLEttXHbNW0EOdhu
RCaXxgWYcb+l9LV29L1AFOPgxno1drXUwDqvdkZx4msE1E46WnBL3PwVW9UevqE6
omlwf3mcL08xbVmFsoiRZDGztVxQkqij5IYD7l6YK3QF6tx8bZd9zGIi9kSfuEEi
QZ66Ruoxjab0nwdp+jXc7FLCt/v/7HxmHuGL6OzrYuGnF79anD1dzhHggMOFNikc
E3PEkF5d0K0PB6DCW0pv/ivVpikdZi86eI44g/0oXpt6feUEYwG18K5tE2acWmwp
RlSZvSd7OkRczmEG2Ijj/FEakqE6jagpFgUDiYWe/GQhzHv44GlytXZIbcrnjPvT
ny0dqbWUpzb3hdvmyAASK655f25SYfgL/bMM0ZUbfAbaIxTorKuEDpEWIrZrxv9V
Grv8sJMdcULUTDY9+eo2iKa7APU5++P68EtEFWEqv205yNuzAl8Ej17NxzFSaCwF
dWE96FmDpMsL8SQBGjlei5Q4SX1P5T7F3jhWuyGQxo8lYBpz7bz/MC/+0rCOZvJD
AQsa1ntDtC54vnTs45saItxREPcwPN0AA20nab9uSTLtpgqLnmIogL3qdY+EQ7Yv
cU1qSdg+fDjHGPO4mbjB7hjxUjZq3Dd90mU7Donddaig6HtPQkA5wUOr+xNlKlU0
+bfH8l/f8w4V/sy5bGjj7VaE5crogUP/5y4LWtuXOWEu7M374vPUOMBjYuV9iSpk
k6GWYjHoFKSgc6aVBFZjp/njcHVQUXa2iqxZQvcMq+AkcUlbmcCJvw9f/pSkikbX
7gpiyjwJG7LsG8aJZjL6kGc3rb+mZWSzRkh8FFqw8fIaNEy2Bs/GE2/CY9XcfkWI
WNNLk8qqoOIjvNwOQ8lgtRwg9JvIVZIF/eTX1U3rWHfApNptYiM7x2jqLi+LU8GC
nDlf01JPTl+Dd0aZxDrMoWfwg0kRdIMSoyzQ35UPX3EkuED2VMmTzMjc8CjHbVKO
uFdOodCvqkSAJuvIynhVi9cm80yz1HUPuQ2XZKIooTGjqbT563Zp2Vk04K1DtifU
bSvt0S+jkDBXPxgMyL56AO03acwAxhJ9COnlUQazleoGv2QLOLyix7bE+Qh87u0U
DumwdCw7FoM98FT0OwS6n/FUZCcNh12FtoDGt3sUC9wlbh1j6NIDkfvbAJnF/McC
5L8kImmtzgV9WsOBk5L67QthTB5yGyAETHm8RB/IoUW3jxvh1BxwBG2enOFUr6be
uTKlBJQyMFKGPtzOiOZsgBo/CckM9Z/Pcwg3NF7dMcMpCurIABITHLRA1JXN98L8
`protect END_PROTECTED
