`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sIFbzdbAC3yfX+Wizlthq65a6DJU8eQuWs/N4GmC0y3Rkss8msn/1Hf9v+Tb7P1a
MIopA0asnRL2cujwmwtq7dOGw8aj+p0H2YYxzwSB0FXrPydZPbC7UOARndGAP07k
5Zf7P/ils9U1Z4jSySPtucEmLMsu2JEFsIcGkO3VikJUklKgzuSHIaCFcUaoEDCD
nixn5gdOwAGBilXpjDuac9g5NDzi6hvcyPM/68Kqaf0bvn6S5trHIy+fBBXRNeBK
RaPtKBtzsVhKchOVr0f004/JSn74IWlTic13v+Py8q/sh5Wcrr990mqD2hrvThWD
hgjYoiv+uR51kCBaDe3bUf4e/SlxqgHAiL7Ok8CxI4IaT0qE2dHWb6RskiP7qP3s
on4q0AW2nnHoSXv2KxV86ykTFlQPPzOzYai7qDLv6kWUQrsxfA46Lb2GkM5EPXe1
AVSpay5uOA4QynBibdi6IrpF9MX4a9Mehiu5pwlvjUyqUdS18iNYgTGrQmZP2bPP
GTW3+YOkYk4ZLNq05/d28Imgr3wnWsJ4xOZQTfzfV1U9o++NFYEzSJfhishkfYy4
lC7u0shCn+7W9r9AJY4wcWC0IFMIs6oX72nWwH5C4qZ9kLvk65HIxkK/DPORLJOJ
5v+naE7rWytCC8a3daghdnvLOLb0Zu3+RHfevTomUnmIvknlMHO3LWpM+W++QSAt
c+XNshBPzMvy8pMO8hY0gbhzDtA/D4ZDtXLglKI6psc=
`protect END_PROTECTED
