`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xelz4nVi4+JXHWztPoGrViX6cmI+MDiEuAWGaJA9dGIu+H5f5MgUkZZgTscsXiOE
PrsR5afBdkk4NQ60CIgW6YOxjcjJOkTUpC4kNU0BRh7DdfLKGUl8wAXe/1Yqip6C
Ph59RjEt7YRNzjXnuNvqERawjGSpT3E+brBrPSFVZsNDNJ3jFJ47ndcFdjqiDro6
8obljprFDaN0R2+vhgNxOYtR2msLrjkJz5IM75MI3drTCeNczhel8t0rnk4CMSwA
xn+LRxKf5a5039KVD/i/fWX7pNOQB44SFD6VppV1k//xowsbzt1K5K/SlJuCtxpK
VtwlymNVSXyrAL1dQNyyHBh71ZkQdOSjpNFnACH2x/ANdogmjK58O17Eh0p5hVoB
JT83Dbin0tFt28loyHfbP3e9T37EywX56XLtii6czJ1p/dJQ3RjlUkPNAIXbFIoo
pxmfeiPMDMqAzWOKgxM5DumGfuJMNekF0x070uBOek8NAfeR1f0u6eXbmzttT3Wc
XG9uE79bcdDnFMX72vjIr3tPQrpS+BcWvJvt3680MR+QCJESp9xtle2p76mC5rUw
z7Qy+261KpYkMz7Ckp5YVlK5X/QlYA1v20IEAd2t/eAGKjz0E+6E7lxRoIVuPk+b
D11xf5mLWVHYnCpgYgymfpOx5Enm3zaepyqzcNpkPNdw77SbpZKncrdmd6cmwWlR
IcDzvBXxA4dP6iB2/Ttn3sCD5ZLYu/Wg0RCp9Os3J8EOCx89RbpE+gybGcCUGVaK
8XvBvzgdXtikkQvxPTN5x4N1BecLdtWaj0RRzL1TakXU9HfiubnFk7RR74iRVoWg
84yOuc8Nzwk9/PkJZ8r0V77L5Dwfk7eqkQ9kkzOn7tohYw6T0GPyauYcOtOeP7Hg
04qEH5OAMvmr2Ce8shuA0YEguxAdyY5nKRVSCjfpV8vMmHoXpdI6jIoMGmgRiVAQ
mID+wmjA7bQ4bv/ryN+tCrH7/4kr+OD9voUYPXntJSRtQpXAf9acTqIT5nb2OhA9
sEYbO1A8HcnhZN67s+qvSag8lkJpbt51Psw2MmQoIGtDe8Ql3pUmZuSdvHXj1ipM
2uLfb/0ZupyOhhsNOF4x9Nw2SZh9BedfvquWSyk0u2fkDg1GGytDFm1E771pMlw5
jo1h3Vp9+eVN+2NqC2OMtH196oUTrkeJnA1TVx3I3jGZbMabJGqwaOsUGGU0VDEa
rdjW3er2pxYIFsLyBCce2pPss4KNGf1m97rOCeid4m840VzVXH/xv9+bNqUgt3xx
ragj7vCVskcYSZI5/a4+No64P1/3eY53/RX87sxTl0s2A2R2KdknOwz8WUVsj0yW
iLrrd1mp0KLMSOvlCiR0FtX+IbafS+j/4OPjJkemB2OGsBPdWjK0hwwgPGLp54hf
0scZNfJMcxVO8No0hbZ3PE5KatdpPd+hqReVeZYdrhUUH0/Cq3JX1t9xFtrAU7N8
BAhW1Oa3w6u+qXdvwAYbe7K/T738o+DrCX3w4a3H1NvVMf5VMT1P50WcKdR+qgV1
zRdWteyHERImIWkddh1NRsHzi4guXIYAj/ql85kGrbD3svwOIkIUiiB2ExYibVZN
6bEzocRhvVhOOQxgRNv2pzQQqi0kKM9DyXjOcS33JPhLdSMvtiqQBcfQ4KTmO4VG
DX+cUyKHkJ6xGytkK4ohRdbURJNXAsYS9L2EaveUFaXy/eA2KVnpYYoRenJi0ZcW
uGRl3T1peZY6ibNoVNZvtQuFHERr/oQ2bLfgYyG4u2KdgGA69atX1CAiZ1OHk5C9
Gf0VTBJ+E1s2nn+Hpgoot7h2bQRjDdnVZRZWbaTkcAGvJSzrdXTNpIu3t08jHJ/1
2dd7P3rMAuwX0eFboVgsD48oJY1uMHMRe9zuFqxMsRx7hA1Uw1z06fqAn0p0XsMu
jYeKoMnW0IzeQFJ+t/1RyWawtmDRv7gRk0Nj9wTlhmf1cKQ4S74Uka4LResoOzWf
g90dlAGMlNA3ErGEvJfJxIZjwa3ffwlpktE0KtRfPSc6YlaBR527wO3PXxZ1oHx8
CKdmFZ7b4UTLTqjeWCczfHtyClOD9LwKnldjmnbnIa0wnK5bya2Y9ihTUgDu/wjj
VK8hmKGhAtV8kk20XNr4ivcqAOG6/lezbrB8AEn0zRgjKTvVz+tGImbdd34ChkOi
xDjW7nmlj7uEe2zGw6KbK1q3dhqzQAf5r2Hq92ckQlk8CLA85D/9lg20N41VOV6N
cLEsAkiVTSyhB9Fz/e1SD802iZ13eEgmhcnEh2WxN0QZ8vKRfDC3u9jlPJvCV2d6
v6BFOVHpwxmUBkCMshPltoAtg6I67MjumvdV98+pNHgowIbr/IIG22RnC+qxc8JQ
GycodsfH+fgMSyVxmTC0AlnI3Bog0AQKGcsb7SYWSs/wwYJbygIengHQEN6OKvZh
of8n75RGnA8E3syMVHgpKvjU9VHREGEiOmDGNPNRZPMP+YmCOUVAeqOQHcVPZo1H
VkXEEVGJWgrEIJklMl2vfO4XAjyNBSHe8wxvCBMsPa9+6K1WCwr0d0lqaarwRvw0
93DUWY8rQ0eh5oJiKkfwdJr2k7AwZFwsBVykwERHoPD+K5Q44A3Eh6ASuF/Qlpzu
jMvXaGkHAfTsq2jNOkv1zAW/K2IlwRzRwQAuvYAxPC2BAvPH41odzRFOE4FS1rf8
YNguf2ODp2lFrS2pAkY6sgP1zyI38Q3X+q9IW6ZQ6fgAUKMM7ezw7QGDPeZ2Cqv7
gqkmdEwGS+tXzRujIqoLn5OSskEeVELt25nzPZB+O38ZeWLajlPCCJVgLNlVQres
IoRybrfChDX4Tb9xrMqV1F5GQCJfOOgbBYBRxIz8OUfCLl/MfO0IK88x4L08xPas
NsVwW8yNj3d+zdBH1EktSmKcV4ned57XP7f3VhbfbRIyjMZTqbsa2tNZTVxulU0Y
htPR6EATj1iKzCMrLJqGeBz1SA9Dy/zdMyq6xB+u994Q47Ih+9DEYVEvD4VT1MQc
CEYXCLeSloSaOxiXLIDEHVT7ZIsHPmgDzI2lQQcmKjzSyvSXL5di6/Pp3HtbkXSV
vMM3rWvPUxqrrUJRyjvjNQCXmqyIktFZmNirorvgB+rO9zaQkQclJReH3QxB7zyJ
5S+dDypCwZ8oOPLhcuTLof18GqCLBStKsMnroTWc4qLZomvZC2a+kh1DEZ7mGtzX
68NJLJy9J06hZ2Z3R7P5TJxUJbKwjp//F44tfCFIktl+OeTTbWdqAMjvnX3XON6h
3/C4S/V/s5/nbbj+UQAotmXdnyu3glLeCIeT3xa6C+PLNLqO/Bwssvw3XyY8xSN6
HSVaao47WApIfXEjjZdwugg/xGz7gO0AE7fN3gWEYTLfGvxinglGwfw3h98U7Q0m
Ni9znaEzseZAQrRnvRr5XHS+BTZpkQTo92nGzuyFz8Lbvp2brc/G+qdaKekpCPFd
vG0O41SJnbgAImwQhTf4ekD6SFBc7CgCn739LthUYJim4CNKDHJ7JwnNVFs/hkDJ
A0MTr5EpCBs8d0k+94jQlj3L5sO6kW1kUZ9Ll3QR9xbTWFcGePpYzNddepS3xqtB
Su3tTtL7jH28in6tN7fG0E8l0Ej7P9POphr9HNL5ADz1vWkn08pjypsKKXf1qGMm
VqyQ3c7aQ1zb7hQxkBZkefzhZEHBk6YBj6TL1HsZNlbCKW1EAEcET71wF5EzHm5u
bw87GJVi6UQQP0cTaee5aq738xqpOnpZZwiLC/RhwZweLCHLIhbQsdGJNsAE0J/i
k8uQlU3qzPHLLPNoVYQjU/LDhc2gImkaxqoTa/JfvOHNi4GDKzxS+MmZ2PTyfNfa
mK6h0SpjACSGB4fSa/MbI/k5uawd7lKPeedWqOfvaB2Iujj/dWWMha+iIWIvIAPq
o7GlHys7rN45LWcBBRk+tjH4rTnKo6zdZ5DTpHQCkslE2jlItme0gZbu7sVNLZnU
sDAC/NrJi6R0wHf5iOiZXd0QfXQJX/yCV7RrRdBxt0Ezamw534pR29WOS/8rap4i
+RdA1goK2A7eQjgy1gvYm865wntQ0RIINlgcrrn3g7onjOh5Yhq+eL8jTMgc/njI
gj4meNfvgBHaTVH1AzorE06vVBqFW0h5yd1yP0MahcrWLo1qGYeEwpPeb9J5Jvt5
VeAv4SCdROXGuXV6gfcJuGCYwPeEvJW+J+TvtZfK/cbDg6AaUTQVQp2pYq1GBnC4
7RUDjAexe0FBfUMVjmxxoLnn82obXdoqArEE1ZHxvP1AJzVNHVt9SNLJweAC9TLR
/5jHCjLVMs0/m1OFe3yUmz0d3Q+OYI5cgprXeQwU1iXXxK9tF/DcnUAvFYmceD6c
qBckR8xEEUhY2cfphslTP4uEniuNH2nkTWSQ+NS/MGlqCI1tPo0pxaDhRw07ZqFo
+xjIdHFnl4qySZFs/bgkwVvsVWLR7ND3nj4Qisb20WfZy8L5a4pjv1fyNO99+Zj5
7uhWWXtm6GOptoCo9AucJ+Lj+kOgDQO+2DwBdboP+fSb9a9uzR7X/gRpKtOR+qmo
UTJ6yWer15FVyrWsILaw+NwAauPwXo9v/Hlil7HAmnOgeUZgSMLmJWfqkqZMsI1L
HK/h/AEpCwzXK1fHtUh6XKrStiB+D6WH9YLC9x4raq3Ev5s0FH+fOtCxV+0fnBbq
8hNFsKEw6bzkjmziUtRahGP6RdHhT9qytq5vh7ZoB6TDxyggQY+yjLuruC4r4HeK
kGcJLN9C5d2mNpNayWs3+/E0CTW/VQbPSnb1Ggv+wmVWEJaPWXzfl4pegsFx3E8N
Cx0/cOBnkssKopnXeK/Isouu8houiOb4gyG8gBdyN+iNVnJNOLpR9uIEnEr/3TsD
U7qH+WWFy2wcQPyP082mqRG8bji7S1yxkhSvuzOpIYnzX7HREvJO5FtiWSf9sFiZ
KrCmNmbbu1pBivcxeCi1P4e9qe31dwdUQ/jqdD3FNlyBNE3szR86RBcUPjQuRqjq
U45jiCiCFFXg8V5XqFQZIUT9hhsYLNFzOyrlJE+SnflFeqaU599GKDDhtjZNnjmz
anMZBjIf6THPm5QFrp32i6H8OxDoB/9Isu8NCL6PHDbY59h5QqjnuZTEMqksCsYS
ez20QqxoAzqgDoyXmge/Z2ORTJncZjAiZidOwj1P2k8B/Lw40RzU9/cuzNXic9OY
ANtKJQxlkNiSDaROrCSOY5+XP5c1eeOkHcFHUDyGThvYWh4m4qyWmdCGd2RSyOJO
9zKURN9czMu0z3fyE6bohdMTlrTEKD9z3x6UMtRa1QRT71mkOmkjEIiq0pC6hGpt
WRVlwhhFNPa+RDMvnvxxV6h9DmyxHw8/r4hwM9gcDRGRpttOKq6DnuMYSzKhtt0u
Y44ykaRx77wH8+OYgFxEJi0krs4UQajRqi+7dtgLAXKJgZP7c3lWBau3KIKnNPBF
icpcKJzm69qXbazJdGxtukk8iBOmCUnhLl0VQdM+t52HoMKiU+wkLeP+k4+8x3Wt
VTixdV3eSEs7JXvGOvpJ8AXs65Kw6+4Z+ail/b7gdOU1CDeqlV+zrbbnsEWQCovd
lpRYGFPux+iOwcVWs+MCrMmBNPCByXt5jDikdkZekpQ7FU4ADt5l+tid8BHv6hC/
9JS1JqX17bWBbpQbl1E7XgSh5ZkPpgo5UT78Po7qEvahjpHD7/mmHx498BlU/kLQ
`protect END_PROTECTED
