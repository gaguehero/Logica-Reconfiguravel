`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPdLFkpOe0TxPZyG2BDd+bfRTuFNN3YJQdRbGTVVN6zVewgeB7kdrl19g8YVsh2u
l8eyat+IWjRw2n4NvJJfzjbkircD8mQ953e9Q4yZ94T+qPukXn3lccpFCHuDXgS9
fvtz2mogrzEfLAGp8jvWJ9oz3re1h29rJl9AApAM2z7B1rQVmP0ANOUsnINxZmHD
VzpRXRDNMaK2c7jmODDqjEOSKdYrDSJdp2tzuttFDhedngnU+Sukjns+OuKtoGOj
C9pi4Cvoa69TccUeKRSA9m/4tg2JJBM7tT29fZktYzFTfoa36uch3zzIWHHXcb6p
Vaf6e/sbX1rk3Tw9/NcMDuIEko7dizYpYMAf4dU3j8XxGaT4akEGo5zk8XxHI4Pm
cHeMPFWLd/oTPlBrBhVHMvGFkmujaFsoU1jcaTj5j3NoCSvjvoGNSKUCWrTKu7ud
I0YEkFnS+fTCtXR5RhIBbQ087zrrV4wbvMwJak18l2tiO2SM0b5KXC3/myzFGmqD
Yo8CZN5in2jE0cSd6//QyYxAGp4igxbgvHSbvbIACYsDOCgG/ushaASaTz7xMh00
KDf2JNguJOOtJ2tFjvz0A7xz94Z1SDSgKHjvlUCHHf5oTDLTAV1rGh4S5fWpmI9R
MdNSjxVdWxeqqke2r9FlLAJ2109KCTVg3sMjKH0KQnA4OkjMUNZ+qcNOkYyLEmZ0
K3AG6541VR4Lq/geWbo+9tScbubDLWHSiH02Y21ZwVXz+YAjuY+SrOvsC2zUtR2W
hqo1GMAhm2dp5rmeq1y8L8cjLamqyOAzsvhS0foJTPdLQgp8nWkEBp8pHlOzpbhF
/uz1sUQZXL7BkyiuYjNEl6ogzWolCI7sxYu/3KFEOy+MqjGv/enTETGf4eU/6uVg
fhxTcZ02CZAmw6XTzKIujn3UfyF84H7dlUCbrLRhgXsXU8kSMwiqoEZl3P7S73S5
4B0KHrlyDlNq0Ew2XB2QhWa4x/oAJYMYhutFzmhwtLY4w/mvvz21C84yW+U2ime9
sCcrTfy8qKVw4pTJDnVWHjCP3/CG4/UC7SeuU6SHQD7iHKApuMzoq3Eh4TCFtHQS
QmQ4M67VOtwiImaQEaj8J+hVXlHY79cvn51yKftYPJHzrKAEK8SZBgsWyu4GgZTe
Xv0uU5PNfT/tBP9f/gEVjkAf3hE5zNaNwCprLUEKv9tmZmcwmJabn8D5i/OE+5hn
1ivQTO5gjrJsMhp108P3zD8wSLuPUUt86dgHxe/o3hA/nlxD5nQMwUdk3jtxl8D1
i+CN0yji6428sV9I2vSr+/Ob31pl/4Nb/rQ6naCn9GDCsZHopDpx21qhkEQlWu89
QKiNeLqPF3CbSyYJ+CIWNRVcrokfZJTS4kOc7h/Gr+buRjL4d4IWKKAJ0pUN7BfP
k5E+YCKc9aFpwUcOKVIrw2CRu36wkoZZGugRRskeKvGoXE1vN58yFOMrVllM8DnH
ufmOQIJ4gfrd7LP/jAaH/gU/l6eMJRBN6AuzhCbfFIbgvSmLHNe4knxlQcRn7boM
FPPnPjbNLqwofHfqKpHPCMZNdN8rIEZThTXGpAunuG/gWbkvVckcEvdQQnWZWPsL
5hyi6FhAUG/xT3EdgCin3JzqC8etuEWiW776tINPf8GVSRgdCsXyBb3V4eCYV+WZ
lNk6f1+3v0kyfkKcHmwh2xWiRz7LaJYMpINflUk/RRqWIplbqLcToc6DMDT5MZtc
cIzK9dDaVwJlbxgpfz0AvrJvKe0MN7g7S9Pp4T51uj2M5spfIvyuQzleu32PjtfQ
n/JFYSR89A+N052qbA4cVyzw3ulrFd+hw/HHMXEZd2neOoaqbDuy5123G6dpDqyu
KG9Gq6Px+VOxJAdYj/79tw/nF0gdGKaou5nvKxgGlPKgdw1wXFGMOlMF3BgblJQx
j4aSrrAi90Nq9ZQGJJh5cu8Ww3uB6jKxifBKkLFMmfbunXyBiWI2jomHVRNuxNQa
t+X/XpCDT22akdMMruslBXEwGHphhYIlfNpH/1qyAG25YSgReWjL6btanFCVpwZg
6/V9McapPgauqW6nY4PUy6yb1Iv4RlNJpKBpWl5v9qN4bYaGAfqDZ+x0mn1WqMX9
e6HOTrpr80la7v9Bw8SMmuj2Iv0vu/TLApYT9k0in49ESd3b7+rdRixsb++1oXOa
ZuNNxf1gw15qJ81d+spwlVY99bpTPmXo1PIjxLskbGP5W6XJS1DZ2mr0+ev3WpsY
b6theemKQylmUTtwg6MiZpHxBOLL3Ji/QFw/eaMz+I3B1aue0G+s1iau30DAbCti
3vA80eEGI7DxLfauYi+c8zoEYiovK4w/5/YQq4cvIHdQR179EzUNP0j2igSV+fdz
ztt05eQ1Ok9vk8192sGg+/SXaYT2kiJ9qjlI6uynQx+w+jKHJCD4U8wWSNEVS2g6
1tSwzs2EvZyKps8Hz1cXKTvjlsedc40gVq98M0u5RDdgK7GHxfWeJfLhvV7isjDV
X4PmN4+s6Vqf4n+W/ttbXbwxVMKm41RrqzVLAHg+Gdf6Lgo8GaUFG6rZPeNlTRex
h28I4pLPyRRss9e3bwZboYgURhrumGON37PSrQcHlPkYr+LkA1cqgRF7KUr0OIHf
eyc29MJFVdm+nV8TMjRA0HOJBs826E01SzgKZrUnCCgbJVk3IBfH14ABmqqjmr6b
VkGYyoLKeDPZskZ4t88A0iqPhPYhuQggJLYRrJ9tcyS+DR+RiGobLH9vOtN3nYya
44UfjXFDS5/t5vTbXD8880kuR7sULrWmROewiMy/oQwha90sg7146ZV880tqaBvE
PpWg6iajhEzZOxb6XuqQtUgAD+gqMJfVtaxxRvQh9whCorY/UxdE4IoLz+OS+knD
DWv9zWnBziXsj3Qqryi0itrS8vX0IWUZLrtKqm/r6Uz6kIbL5jBajJcFM6efVJ7C
vz6QfixXzXQaocLVZV15czxaBRxw315c6kv3VtKmRBT0jg2yt0BRSeSM1wBjIWqT
O+AHYrOfkvbBGZ9vayPmS2ySA+IVuOtklwAi0hfb5I8CFw45426l4JB5vN/dDCq0
oDwSw/RAyGDTrP2gDcIa3Q0IQpb/86V7EM4cTyoDZXw4t/wxHfgxhS6HZc8udnw8
09kHuBsA/mf867NwsOmb0cl+0BfCybxmLk7MUE4q+E5QfV/dTHF0ZXJud9V2fBsy
xu6zTA6MOg25YgOkHx1d/zloK/Nk0J6M1d3gnpmr/KBp1FeZO/BACp767Ec1vaA7
IcvK8YgxYMEyy13Gi3S6JEfEvRHM9CiM/67vth4ioF3cB0qhFQLOosT5emN8zofS
fIr/Fk65Jwet700OHk2pTa4SX39n24hM2SHdOZBWuloUT0kGGMf2OUN9bBXqWbKQ
PmIcymc9dbDKFUKrJU0SG/vRwc2MtIaSDGlAfI7rMu+u9z/ZiMPgEC8p5k9zt5k1
mytfLIrroEPsnZTvcfW0phxuq2UKX4FzDDg3oHWlvT5muGgxSzumN1ML/+6VkEM5
4PZMXtNvuBvPkWAwzBG1QOAgGrAZH9Jge2rBvSHw8jiXS0nC+8bHFqoVkArQJw32
RiVAMIPwq4hkB+s0DD6Dx1gqAEgP12S1rWBMVnd9YRe3G/NxvUKrinjVdl0a+FRv
Mluinm9XR0QEWvTMaoeG+L5c506x/LcKIVecWRjvT6ldsTNxqj23+zNE6xlCB+aV
UUdPV88Fpk20TS6srLdyfttfIWh96iHjxVbnbTby1zfwx3s4gRL/5kPGjaZtRA6I
2Aqyfzh2gyQtEJtNq/HtvR8+w/ng1GUq8jkkDPFQ7cbYgSsFhew/4kRoh1UWXZYS
zOffV2wv+RCII1X7cbETvr7TziK74QRyPK7K8lf7nOt72UgR/YE28ktIV3MGfcjH
HuLEMv0B77dcZYol9s2YAnQFf+ggZTc62QF6lVjAiqiVvYVwDkMqaBk6aN+nNlAn
knuHerKFbkLZM/RWs1HqDM30xxMvCgr+CH8nT9tNEOJ4ML/ZdiRIP5CYDmH7+19/
9VBFD66gHqN4RjsP8aRNHmGtpL4ufrcMjZNXh/3aEx5afkl1Eh+Uh96lAVOTx+0h
FGX+ETDxn9JPzEkNCJCYjBbW0rf+thIWkj0P7arbU3peQ5ckpzpE4trNWlB795xc
Jz5Pe/Vlu5ZV2y8d3d16X9vW7RQopgCDXcJh0b90C26cxO4C0DDlzqMUdEM99sdi
bW5Se5N4JAM//7L7LjOBk5dPAMAijIe9f0sBqQz0esBcLV3O77W/5VxaWm+gpkAQ
x73FHj/X6dNzoKLWDP+Cy1OkViyvyxNQ2QOiX70XHYZAjJilAb0dIQYmMYZsJzvF
A+jJDY6ZGOAHfvlbNS0rjfgOMZZg9Wsu8yBARn0UFespjEelDknUuOmcuPcc031N
/HsEyrtJJxmOVU0rf26HzAaEdV+W2/R4tGOLIM9T7vWqDA0ZGOeWUPjUH28dJMEZ
N7+r887z/dPolp2SILpTMYtPNlCvw1skcMtHroF9RpLPr+ynDy2E6syktQqcj379
uccuxYoDTLx4UdGVL5GQiKkByYVSjsjMA+DEDEf19nS9ZsTMSdUeGmlA8vAd4sDZ
/t7OZWiiCAhZqh9uNrATy1Yjra9j+OFCwtK0WY/efaJsm6wq2Wq9EajZfu1nx75L
4ZDhanhwVNs5jcZ8+PXjgitCRCmzkieSYOkoQYeWODwAuj0/Yq3dduVmpNquQ9IQ
Gs8c/j4arG1UXsUEbpWeSle614xuJ/SxuPOmbVj4hKrnrOYsE9+TJBN/ca1ll87Q
19OekpXJkTQg/nxGU3kpac6XTyR7Uqvw0bZR7wWRiw1EzwoY7IT8BcmI+KZ8uc9D
zh2F/ZGkEG63+R6DR71oAGX1u2JhQZz2H/ogWxcta5m0/omB7n/gqNXQdBn8lgeh
KDVgPn6uENamMytaoA1qrmQJ94dnq0YOLWyZ9huPUVzn+6+UYwh2eud+hC+fwf8T
s6WRs0S+0eIk4bQ7927t572NNKTEwyGgpqe7MJ7H6tX9VFm6t8mFefYQKysDwpJr
ckmJDNcWNH3N8p/A+7zlWUDkL3a/2Nh4ex2zkwTl3Q822csyjppJX6S97QawsxKZ
rkvxAIzdXH3VP/0QmffPWzO6Qn9vy2XavGuj7PrumrR76oPZ2ZV74M+uzyYrLJcM
X494gl7OaIg3x66eUXuTDn6BvicljYloW2bWidhk6eNC+WWhRgb2BDyGsceI6Ijt
NAT8PcMD3FkRJAf/ATsPrCbTQgBLhC6R/6Xd0hIscLmSHEz/HEejb83TwWor3D+w
M5GKzKG9JrvGe1of1qe3dtvfES2mm/vod4CGeL5PmW6ipQApR5Z0XC7VK8UPcV0/
45C+BLpobmeDC3zshoChEMP9LYIMnsL5Hi5MSK1U0JcZOo4AZiwld7IVrjRw3CpG
W7OnetuPKR1GFNfE0PCLsx2TOKiQzwsjndI4O4zuJ5/YWcF/egy1j7SBFkYdTgWw
evcLNptUt3AU/6ull3FlvG3ipq2hActkfzqnvDC2DQE+oi0OQBxpBCq0/8ZcvsL4
s0NvzTDeSbaIlb8Fllmy3/AzxpCjJG59uCXDXA7SMYUTt2neczyvmmvtLW0Egr1I
9FCZkDIMAv9PPFgcgsNy8K1CrQVCdWFF4lYF2N7xnL6rrM9p9WZZ2rpQeRHx6J/b
oGt32P9qA3X7h3QAyd7ibbIZi2qvTOOzo3Z5leevlmude72iHnnVP3pBcH7mAtA5
k3CRDQVknV04f6/HR1VHBwMoeZU+xthkSHTf85z/WjD3eNnDGLlnNAr6SfUNfkzR
cZ5YIIP8XDo3G1IUjfUYXdW85etRQYzCRsQ0EIE4bumKrRt3NvRPZa38H6PKRVtC
52BuUCjkgizlSxrG6ejF6dEt04l4NkpxNQxhPRR6wTL1dm3wtxPpK32/uXnsmVnQ
015PjKfrC3Ucc83FztJtKvce3CSy3Vl98mKQCESdlqvbYxkIumikHHTPqf7MVxfe
kdkAbk7En1NpyvE/3lWAZnzMZqH4jMbgvbRH4icut5P1kdZfQJV9BP7wz3sVcBJm
QdKzOIMCeJXZLBJKjJDZCRsYpve9yJZwCoA63iAQ/OhZO8A3P10p4lu0OJdtjeJN
n9EFk6aQXrPa/ulvnmg0ULxaPLNMv/pCI0vWIWvOY5eVTZSC+QOoJHIAOr+NKB7a
4pGhTcekOGkaCPSd30v+1hOFrRAUWLFRCG3GT593MnuZ/I4akY390WkOUFL28LQ1
BfzUfaJcRhDoAt1/yGWGHY7GKEfY0ebX3pE7uNUuIEVeSxy5i5xi2f/l+NjgXuPQ
Id9t7QykraxvZGKBvvj9NNdEOGM2NzCTfZ10qPrKCr96q95HD3WXeUrUgJ2i6j6R
qUpO9LCPQ4vBrrYNuoOGiT6i0OTF9DFbBbcFc69zJEqJDt9PTtOpKP4OI7Mi0LDM
F5Q014V5Wxb8FPAWx3Fd0K4BQrAiNoX6Ua0o79HSt6cQTJxangQk0p63q1CHMKsc
CEznmj8nsquP7qE7sqIy4AoI062K/gzyUK7n5BS0HiNRU3tKQSTH1/ehBLwOl23e
Y+wwBXFWqcPvgIM7oT+Aj4gY1hi+IbtwkWR8COslD5/PyFz8TCA5zCOijbH9md/r
Zj9q0Rn8ywCScGQAxvuwhBLrfBEqn3F5aHspJAOiWl4=
`protect END_PROTECTED
