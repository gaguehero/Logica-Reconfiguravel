`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LSWb1Fa8OtsxQZMvBbvEUeMOmIAnfPI3NYYE/MFVpAQGJQuaBmtBM3nePap3id6a
WC7LzpLeF5adRV0DajlXcD/aQZ/y5Oe3fAgRgdneTc5YMfIFbcb5Ji08nNJFXvrp
EymXP1NSAzlUvftfYQ2KSy9lirXGXDEpG9mp9Oh2iXHqQ830+T4VRgYfHgIEekdl
TYkUSLjdbHCsko+VI406+qgHWmQFFPHjvw9fw4xApaTZqUlWnPwCu2eklp1v+xVN
wlbWAwRSucabvKt6uCb+y4mMOP0C0WwKJcHDlZJzzly4ADQYSKO5+JrzpZLLF5ah
lzgKbtf2MvAQ011eD/nqZ8V6CKrHVjAEDS1KuomY6PRojY+vmwxpHZgi0qORhanw
4f19Rt4FyVkYgZPwru8+ANB1ZPoeHy/njy25afGXiE+BCBxbYdgLq4Ep3ZLdcAG1
wuxMi3cjFaHoCiTVdBV9HjobU5BU+ee5VwgZCOGlT2thKohMkPcR9fHvJKTDc0nT
gRfYMN2OHveNG644c5Zs7UVlspBEIHkvM108l5DF8IM+/8d7IUxw1Ilks6YCTm/I
MVpJpEnSdmDAJZeUglzqA8/lIayycZhksQSJ1ENyjSLOq5qfITXaOryoAt+uTV2l
694Q4uDkaZS7/RS4gP5SYhZv9qOPCrvNexhIHvYkedrv7BrW01WDvc3rL0Qpb4AM
yStllCAXuVgJ1+H7qewIk+OepgbyCSVcS4cTRrR5PTf8kNfnTmIbj4vcvWIvuDzp
Fmf8V3IRjN2iEZNd1q17BA4ZHJ87Qwx+I1oPh6vYCV8jBlMKMYd2ZaHSBzUPUVCy
4/XGSbuaLvj8ysCSB2HBWPs/sEZuUIdW3zuLYkQ1Su8ScHBLI88md6wWss88LQyl
aExAIHywlbFBHNVIItHPurZDeCNkARG87xbAEJK/sZrutVrleUDf8gAylcD9OO4E
u+JVHXtm5YDIiuI4ZRrA35bIfgngvdVnzxSGM6eQKQn0OgSfEAeX19V5fiZGZHVS
ruuXUK5fKnJDW9Q0ydIkcsi4aWGSDREeTia9JcjUrcNqWxxKawv/bCAEfNp29j4A
1oLGSxa3l725TRsCqjgK+ZiFVabsMEKYU726HYgY1zK6xRLGxhGMmuKm2oweV7rF
L+Nq6y46ZyaQG88xdRHrp0gQGUo57wp4BAZyHCw+QAMGwRuij/erUOdN8TknnmGJ
oyVsHwXjVZOvgxhutO2wFC+IdY+N5sD+t1NRKbSzdiqGJuixf15UhZCDRuCqhQ+J
jhFu/j76JqmQQhWbNCChznH9U4GMJeqeWVDKprxHk7cJeVC3ipmOAAioxm2zVQIk
K+Zdt6L4jAebaktQlpez91r06hyWjgG9RKAfraTJaPmFpsBcfmhRwu01GC4LfGxU
o6bT3tyzlUS1yIVOkPqjzyaQPH8o5gA+jDuSPPkoZU8N7X3cqQpze+EIyvv92nDC
1y6ZTcHUPefhCyuiNBOaeDsovJMScaSfUA4F95K2rbfI1uEnnH7knTNCrp53qlgS
5G1kPIZHNS/O55P/tcA0/ZNXhtZEV86/nAjgP8wNYgMWblvzzpf+n55m5Pku0xfS
gES42BZqfNBHStflwjNuqE6lz5lQ99fNpYflUFGZpWFGAQ1vX4nS+th46O5ahEfM
mUqZGPJRXuBt571uTFjeR68EMowvkwLdOCgRd70cerscRt44otqFc1mr/QcvPyol
fwWKx0gV164u2VH0+041MrAsi85w7wFH7ZgfbbkmsGYoCwt3f8ZfXxwpf8RD2C3c
1BowydIf02MvizVE6zSoQFi/fesiYgjBifCeoaHPmY1bcEgxuJe69Biz7wrjTErZ
+SzBVTnGVyR9+m+9LGl5dxeWfRpeEqsDZNVrOg8DT/8amtTbeBHL3HKQxF8TkZ3H
G2tsiyjvYxQXeCDv/nSAcTNgUV/GkQ2cZIciCJDWhdHKeYStNeK/41mBU8JS2Ayu
JVNaJVOcZ8hG32i/VteN0A==
`protect END_PROTECTED
