`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSzFTTvPnWAjBhESLmBV6yPqJ85htlZix6QgvZTzOOrnzNssuELEKnjmdO4W+ACM
/YIMlQoReWYP70ezPkHm6Pv/mgMRiDuwGu54dwDC6FAOuCqOOV35ds3J41bHX6Lb
IxGIztuTxOJxFm6+ywevAyRkXZzeYKgVib7Dfqvuwpl8xUjcwYN+VQ6A00DzRgso
2hc9VZgTI1eXaBE7w5dt+VPV1gntA3nn/37DzHi58dBmWgg3b85mlmdBstmHKAZY
GZdZ89nDOgv1b+vmTBhWkiOBiFTxgeuZ04Vx7LmhnSybrY217MKI0yH0fESwgQL+
sttehgKZgDUmvbHJMABKGyvOcWh+CUV+nD/fcpXQk5osxYAgWHPjmeRQHqSjVG2N
iekymR0e9kXEhqYoQ+GaxhPr5fEtXK+irK5bx2aedH8cSYXfc90RGlgzFyjj0RHi
qIt+q9e9yu+jw8QKiwzziY5O4rp9T8Hw4mSiPTliR0Y40wSfCU23StlTCsiDoFaj
ztsdP14kNPw/1vwyeja98VyK2/wS+nf4iq7r5iUB6vdYj0uKks1e5jXX0c6aIAZf
l5Tuu3A7eYwW0gVznx4zLte7KkHBV+T1k3CuJqqmTiJPs+grzxhRCyAczNLgR79X
EnyGzY1oI0lnDGddO2od3+uSJuqRFDRIcnEOwZEma3jeOC4bo8f2MTGXCtuTSOrN
Imd/J/FH25cgg0IIBCzK03P5HOg5VG6w7qV5ZBAajogD2x8100f1ElTb/KLJfYYN
6SwvS8fAdS64I1LONxL2+32uu34MQPR7ZIfrHXXMU+e7aRlRpE6nGEIV84yyJNRU
S2yQ05f7/Ol5Ivle9Mcsd54eJvODgnVy1Bn/gnfTSnL7tYluqBWTqu5K6FXKtMqQ
oPo2NnL8Y7mLb/nV1oQEdFO171sEB0NOtNe3lzt2NueMAwkAwh/8Fa07xQIHKj7P
otVIJt7IysbKXABO3HlQEaBCIOhZlkS+ZmyTXOP65bIux8uSSxKtYikNwpsyX/Iy
tcHYE+xPNo5PTtzw8uEUuXM4qCAqPcsujwuptkG7nRalOqkR2VJnx4s/krNdg4EI
mrtZGxW6qrjrztljRHOTwkRKVs7rXDCsVoDSx9j9NLaDkthYm06mXrp06efp7f0T
sLPTRVV+6w4wCjj/m3QnBiDa631JbCZr3gH5xUONvux8KOBP62MvGgKdddLfj89R
fdCOrtlM+piD2gatDIvm+WGb0AsT5AygDZWoaFdtHUgjQSU8nMLNxxM3VNOW2cXI
RoeUk/lLJcmLyvDiDzmR784xQF661N47iLLbZvmWj3PZmo2WuxpEgCJ2iUj/UeD6
ADby8XPdARZDRMGgKGxpgq2bdXCSc4LYygB8T0jgdZ9yziC7oO+MLQhoVNbl/jg2
U+l6+tGinDUi4KIlHzDo7N+ZsIVoWu5T6vWnBuGenm6BcpR7Bih0q9Q94peKvl3p
Uaa8XQ+4fzBo7OT2FXNZ8LCekUpH7vzOz7ea+rIoZ5iY2RJE3eepdKI1RWqNriui
Waz9hOIozT3XVVEE4vN/h8w/FYX6UJlog286BKdVu613UE6MokwZUEn7TUkvda+3
U3JWqF3OiB+NF1xBJz0JlcKmMQBfwHjBztYfkKYK2NQ/tuDmtJqMN4E5VmCgwxBI
4KB4ntLnRlWGSLFQ91qp0JNc6ElgZOji5dpKsULj0BzvTyAcBl39hIrARfaBVQ2M
ITJotjGoFtUzQ5+CNGNi3CvhXFzq/58DOlR91LCtoaU88Du3mi+GTbvdLUwUERFY
xg4iBcQShoEtDwHb1QShH6pj5LTfUAwTcn9ae5J0oDTSukMHopQ4JwGxBTVpjsfg
BmLvr8aeyqFKjK9pUNm4NRKM0BFdzlU/foVRRE4P6KCRA+d7NXtFPZtyZ27CU55O
5HsdxRJFEqBx9BP1FiMdCC+gqyGKOrW/U3Pg/GaXBhVGLgFnUnWisJYMcn+ImHOt
9nbvw7HpOfrsN6aOFHTty4s7o5eLB4PN/bzOsDRNMbwUqnyXeVo67LxC8KqjkaEM
`protect END_PROTECTED
