`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OBm0Es/O84+yCsBthpg2RYj2boMSd7ZPcG8mvKrgvTpUynwoNJtKd7m/3ZbhzebR
hsHb+EQHTbZtpngQnCor2S6P6RFqkJZ0bBclI2nR+R6JDPNs6d35UsXdDyTZDHOu
LxjUZa9ag26HRqJu9CcTLFTFcFxuaxglwoS6+imQYsqIqX3WKU/AbvvZi91Esxwx
gmq/XKJR9uJwQmqKAbrRy430PKMCrauP+CaG3JTEcHtulTT0stLa8X2xeR5vbWob
EBI99dMbbmQJgOTRaU/zNsfKqZ/8AV2bKXd5akvJwLKhm2MH+iJhcRdTjZL19bmR
ijt2duVydsjtLPPHSU0JrrK8mBa/VCEOpEsI8ePgcA7C9RH/e8HVZMSXp2KoiP78
MyG4n2L124x3HFYdTGSvFfiJgbOw693n5Rw0npTrvT2qLHv0luPBIeg7ko5yTXgD
CtrpYgdgZ6k0o6nCClrrmnAeOa0Xaq/XrFaeWwXt/9wTP+RKBk5E/99Ga89Nmt6M
h0kn7SDy8ftcY/PyRUkrEnhd3O6c810zPahWzhdQuQ/gIf9F9MlfDLkmv4HdZeRJ
6Y0KQ0utjb/cxi2lH+RLV4gMO9vI4lyBrI+4dhN5EMPn+5k5GNCMdijy/7sv+4SW
UMjpfEPbl8FshfJqHh7DwDC8tJtu/b/hxwoqq3LfLfBkf9EQ66aZGcsp7a4VpLqn
`protect END_PROTECTED
