`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIO/59duxup9nLXN5qdhpYk6dLhxgWvJc2AWiHikf6ZL6LhY/t9ON6egyku4c7na
v9UrttukBcUgCUjV2YYVvByeScKISLFN8qhiPnq68FNBwHEuw8sV5oJCw3nFdfPt
6HpVy2sk4O228ELh+JSXtQl/LW5rtS/atYqTozewexhw4yUrCtk859KGrX338AgR
qNbCXHuNDMCv5IosLi3e6FhWdLRzVEkFdByyCBIaqxcK0pOumUbh0QEzBiUfX26f
nmb1DnTweb9FEmTK+f4xQPzkIMfo0tNPzRnPRnhL9rmqza6Iso0+jMnzVudQT+/P
N284ScHHvcwSGfuEd0Ws8q4jMvFn6mwFnRPz1HI9Dr7YbFKgNnB0OInm++Y3bKa8
WGQBqZFiWbV5c6w8STeMDLW/Mjq+OiiwzfxqBxqHmJhihymnWZVLMsr0IWkguKIr
mcLkUI8xfrvexen4sbddmXTgG0z/6TF3bzCI6/JDl08Aa2kc6XoOYc9AXUO1GNCn
qKAj4I8tyzJWamXT8W90d0+r+aHSu0MI23muEaBL6J0hd/Ehi22tVvJ+ow8B81WZ
CMtRdAQQC3wk/bzEhKF0vXRpYph44Z1RZioHOhpEx89NY3KZl3oyZ4Pc9Y44GylA
uATYD77v3GNXKjcoVhrKHkgjGgAJIMxWP5j3wu3nv0xwm/lNp0gtA7Et7vRX0+MQ
NSdfLCVHNcRxeowVB6zPLFJAvuG6A452T4wMTRtcYgTn4TaC6Slvl4yRmf/kZl95
NrcrH/NW5dJEPAmKpi6nJM3W+FNTHvGbkp/GTORKgFGTTAJ1tay8IrZn1op1iglw
VjRbT5cumfHPCqAVSyWXo7Zotsc6SDJe3Pn9n07sepCjZ6pW0drOy8nRA16pvqci
pOjifZBqXXxJ6zrcnta74GHtfzvolq8vrA35mLOjDBV6DOL6z5H4bMthFnEsRDSD
9zNBtbvOlEWm8Au+ezRdnGN2PuLrbwoszXWfebQ6ckkj5oh7apMGaNQj6H8obAP+
TOWydkfqsr4rcuwFIozMIE7gb9Gn/edn8ZaR85B6SoUC37Qvg+T3dvd2LRX641sg
zcKtNLhFftwlKElcKKZuzvPLM8FhgnNrdp8eJrBHgsNSlG9b/hIMgNro4hTd+INV
OarqR9AU5Uq66OJYGFdd5Oj4fpGInxo8oTcgAW6ON7A9JaZqKzCl0x60vQOC7jfM
baVuIBTPTKEO19oPYLjByk3DCQUChb2CNz8ChqJg2YR2+0gBnSWY4i3WKRvtxYA4
PL2bK5owg6ekIl4YW2D/Y4t1qud4PpXYDh73W0whsc+Z12/Gph6uDQNfWpyB4VER
yWhQbGj5MOZr9DTotQwpw1AqhMo8cLbWKYz3bx/zKKV8ifUFl9vcXim/GRldmCV1
yDc/xq4rbmWIbLWdtKAvRSsHEgRDqtFKfQvuW2SLsa/G2Cmb+PnxIqg1/aa28ekS
XHS7oavshX7SlP9fkoLTE2Agvxjgf8eJzaNgEsTbV8JH2CRo/5udASMr6wY3Cnya
zKTa/LG/+Dgl+G341mxreHOyBEXZk9EM/N0POlK1QRBG5n0JAImk+5WqM6EWkg9K
WIztInmpJSFukqvHM85sdLNoMtAwg+NhCT8765xLCaOUAecCNjtbLCedTDHyvX8t
yZTng7uZWcq7uxUo6GS2ZWUlng7YIUVOE4GgF3DLuVVlpXzWcrAzhLQcOZWSFqoc
AxeQYy+fj5s+lMx0ivutQsiEmxEoODevXZAO+vrAzR0u8s3uKjUJn5G3hv7ZVx+q
BXCuEw8OlTQRUV8iQ/iuejoTbAvcSDKbIsXR5ykZJ06bXCqwqN4iRCuxEi3RKpV0
uYhcFccBKSAsrNd2P8PDOxtcHhSG5oEPBs5p2ofycqHCE+5fP+YGCZWYlEzCdfzm
YHk3MByYfMioNpnL40uNrumWN5091AcZ9q6lnwiK0yukkPu54kiojMEudV/StSFi
/ql1k84+6mjHZqeXbZ6SuFDlBsjgQnNM0K7R/kMaFyZQ9BHFWuSIy6BJdmKBXEAb
MdqMdbhmOWneoE1AZgMJKZbxMe6dQiq9LLMNLvrK1s/Y2LzMU+HrfyRsiYafI2Pq
jfrnqVamWtZbZrI2vNA2MS16ApWsxSQrG5lXr3M4lpszJXfpSsdR+Grba9SL7R2L
IaL0I/PPTCTnqZo2pIAyCuRjTN6G0Q23FtHexLdjfLtKEkU++fY/xv3dXmQT08ti
aEv6g+VE7YJsU3GoAUCcfxamxrYaz5xe/ZVXs3/+zMP4cbcmCuN5SGsmqy86IPG5
dm639tdiPE+7J9R4SumAtIG+AuGBmilOHHO6WO6Kr/w71p+hTSXbj6jOBIG7XsAl
fBJpvE+77bq4w6UayP8iKkWk7niKszluk/Rx+uOLWfDhiZRTfOcoJElaTiIJdp54
p51MV5yOXvugXcYCe4k+8prjdfwI7o4ki8LqI6ll06dubRH7jnHug/wT2ZjGNCm9
lW2xSTkEyNjJ9TVNQIToMFTwYX4ZkgGL4YxiuSEhY0se7AQNrT2dj0JN44i3qKUa
+3JuVTKkPFhdTmJkfg6TsP4rRpJ1QaPwqYCF5RuS3XZ7vp/9shJmFg13Ry+1p0E5
iTTfZs04CNS7MtoC5fRV/WZYWcY8FElgGUkQ5I2cLK2BMJUOLh7H4mk76YPYpOO+
KIuX9ZE0Rvn29iKGFpYXrpK9wfQgAOyRmwNxk6nGrwSy04EHecnYpUYSSEhb7Fyi
r7cEkvYMhYtTMGKhtlWF92GWjuyER6wPUpObzjlPGOzDBlmOxVBwsRxQwNxZJQdF
uRDxnvIQhykWwWAYNElr7tMMzJEU39VT87zbifGIS/5ZKX4hUz62D7WPArfKH2Eq
HJtYjSyq58AUN7NTYDnJSe5W09ZjfcSYYhKzK+fEtdBpUr12rV/VCWGqeoV9a9qE
EbtQxSSVMFN/oByDniUkjU6H93yP3uUOM+10njivRSlkiGB/2g0uO7tx+rZbHGEm
6sLryuMkm7YfMk/zC1sogAjaJ1+C4cKDDdrFWq62yo4gZc62cVjMwTwEu3RCO9xx
R1oPxnEaspp2KazEPgw7gkhH6Osmx0XL4VmdwhN46h1BpOeJjo81miYZ53NGrNJL
+dSIQ+36DTNRD4nrBNiVRjTLg0WQVlp41A/6Q6b9pPwlgq4aVWFSDoax6SZi748I
0XjCwH/mBY+azJINxXRufTJ2nnDNjOC3cyiMIlx5zRSulk4RwrzdMt7h2C+0Dm7U
KS77XfhhOf24Z4xOaNOywjbWNqmGBwHtlR3LXx/1DRxbYEDgqft0meVFnMR1OV37
r75W8rYRTnP+qHK0EBgw282kDbZcUWQp5P2GEY72spWRYUvk4n7M/qKKLKcpxH5L
ikrytMk5uGSV8fnXPnEcRcfm8WGUUvCePHp+A80BOIxOR/TZXgdm+NZzBsDSXVZw
kGMg+x/E8grD0Y7U+lCVMgNJoFPFtattoaqgTr7pooinBtX6olqCyYOqcnrlIhRf
PHuAQGZVaKd6nw/Xue+oFEA1tUy0R+wAjEyiYlEEVB8kuQVbk7Ttig7rABEdc/Vu
iv2G7EZ4BHR0Cd4AO2UbhcXXIk8qypt95sP+VCz8cL1ItrDY5Gatq2YinoRy1sbh
8rYdtGZuX3CxyqywHqIkgJK9qJkRvDF8c/e4n5zjmWhumdZRliRrNYJM9y//mNyj
THHNY25ijyOw/BSnf23HuYFIPoqBXX70TKD7kCDfp8Skx81BhKBRxLeKvb0BKOvt
Uh7cfj3cp9NiueSD++ItlWgYucQsu1MqJqkDzcORBkSuBl8RVSv+0liMdvQtmO2s
yXoTjT7tC3FTS+0g9FFrB6nfQReRfwAZtn6d79gvRbnsDhEggphKCeAXFJ17y2PG
YeSoH7yy/jYRZxzbw7nemLAvEFMCPQTuQFROTaVIApTFJRG2nZ/5iIr1dr1KxR4N
qBYsiSbnNSqVnJwVR5Qmy8jMKAV82fJRBumN70LjUoXJ7TnzWtny8LtmtNBbfplF
KXwbC4GDy/tppNS5EDSRR/ibsR6vrzlekbgY6PObmwcQ70nqci2fTwYEZ3WKDQKy
6EaFHtrCvwmvxzQKPNSTNMGJ45Cr9nu7ZbEfi0rqGpnJywcLpxI4uu/VPGHEdUgi
5hEsVdHBY3xL3k1G2FOIcC37I6chd48ppuEZ8UFfA3QQiddZ9dwscoY/5eYuhzch
owCEWn1YaIZsfKmK0SUb4yJqlXrWVObq2Ydmkn21BzFbMVtAngowzxM8NvDPhUh+
ruKmlx3qve3z8swUCX4qKvf13OygC1RjG/4yToqEah8azJiOEM+uh41CyM3vOgO5
P7A3lxur4vSZo1LtdMuExC9atL4euVlNnJeYItB1MisotQDxyDqM0n7dW5Fe66GP
W9TqsNNKgtBh9Sjs8nfe5E/UqLluOres0dLoIsua9q+StSYEe2gZB0flfhkyi280
jK30qGXoFb1iAniVEMT6wGDAMTI3IcjZkEJp+171HPfk+Na31i7/D6msXjo6ITYK
gbYgYlMa5j5Zd6YFiMjrhm4gDRQM5wg8kuo5i426WCvfB0tAsJJBNrgE55guWP0z
HTcC2W6xrhcX+m114XMfJvGhP1T8SrNCUUVmdv3agMyscBFe0HvHgtqISvcQLZLZ
HSZa7cwQX9yjFWvebLMgIWF2xDIKOr4q7U3B9xx+KjmycAKQAio3pLEV0c0F8OIk
EL0xdynXK5zIW7zJX9C8sFFvIJ1cSlCo2dSZmxBo4otp6l98E9OW03gb7w94xDuE
W1Zl3BD/7jWbGMwCVWH1OpOfh3u36GGkjeghGev943YZKxtOD7HvZck/9adBPFMe
or8PYJ7bXXvwJPem667D3XLNAM0bHuGZSyeuJEuHVhOexRzYTwr4B42gyrxR8cJ3
ox/WqwZRHBT88yBjAVEfIUuaV2+PnKcKd02niCMqmzrl+AgfwcfODMC5+wdDfiV9
CwXas8S7CtXbJiW8b2r3tJG8NQUW/7yRNwB9WeDGMh3Hpg/Ge0thWMwy3toEWEOf
RbCl/sVBOUTVfD4G4tQQk7XTlnsiZzM6FTqNVgnhh3WXv3y3qZduWnsWu69Zc/Nt
2dXGvLNA857m3jCFlei2tSlswoC5WdmK23e1VnDVlw5Jq9KVLqyQ4tFcES+cZrcg
8eEYtQ2/R3eDZ+QF9vcplqShnWOhYku1EZPZhzJW9yRJfCZFeyJSMlJz1N7tBtnA
G2NyrpXCf0XQvo2q3aNpsNLpgql56Pg+mtSKqIBhfDZOc1Tc6OUd00Fx3HDRqJmE
eRy+7F+otLyAj5RwFfysyswh7xYMtOj2IBduY6z6Yzhx0aId1ja3ZkIuzoRvlRm2
/HBryj/vp4watZq/XBLulrtknS0oBRUoZzLVtUbSjjgntEXLiDGzFAGQLRegxegh
BlF1eOKKLqRbFqXVWwVR0GH742gsEcdJRmKNoMAns/Yvh1Zy4tfWkKA3kbOH+CYu
N1Nz3hAYsX63Cc63/tc+iMwlIrdNbwbPb/be2dqkN6ukzNH7k3+GER22DyYmvwbi
At+2spQmhNNJqJ+BsrjCLUlvtX1czm/klA2GkzP8lIBSoPBBRfTDycyCLFc9AdAv
OToH/B/B+7af0gxl9uwqfZoB0L1Bb1G/Ead/TCWz5DMtUac/TYuB7XoQhdcGPYrk
d0NNdm3bcuYG+8v7tq7aOe6IgAGaDHeFlc0XQd11pi9vGPsH2uu+bFJR/CAF9KQK
opXW/lA3CEqPzMstExMKu2TFIVDrAKa34SZj3ia0KlqB1asPc1kM5GHGTSZAgt2L
b3VeiWEdXFTtYHFIoI59pNqCTQotxzkxSCi48LlTbAjI4fxGcMsgUFbKRAyaZw35
AH+b/caETXUHeV7rHqhNtYMd6aLFxghFugWFXYndIDhD9NILNhfB8DjTKOOAoyDz
7hPUpDNC7TBLCdr9r1Wzi/mPxHUk7MzVLsmfasnUGw/JSJjBrGDHrkJRZWIgeWj/
gNGh3SAGIW/Kdil/aF4KFOn/J2gYPyJjwEelqghPF1/3beZbaZ9n2vRiiMKjOpZr
8B6xp5jtlMkkBoYFEsILqBzTSGsPwHXVzqYjfT7SOfzV83LRn96dsi6M9WMJmUD9
ghINCqbYHOX4Y8fvQOWUtxX+EXTrQJO4zOJYwVX11EGQ6Zn506t87QVODxrFvs7e
t4Vp/bP3/7KcTm0HGCkFPI7mo/7aR3ldewLuYLkHM5bu1LzSKVOSImhZTZ/R+B1I
Cdd9om5PqMaDj4hoqu02tAD+hO+GFhTcGVVImjxnC/W+KengiksfHD6CDkw+TWht
cKdpy6mekP/xjnHRwj+XSDlnwF0tqLwyQ+KR/lgIcKG3uPIxUO/tzxIzQSxqCB2r
Q0cJlx0a5AQaX//9P5UKYOtYWNgl/7kXPs2ogmvegc3Ssp1Lm/eIS2ZfnGTGvXVa
nPGX4Mz5RhnVg6lZJb/F6aHCH5djghzkyf9ozy4Up4JBML2H7ZlfH6AoLg400C20
Xa7HmyFflPov+i/2Oeze/UzbIJZUO9gP0RmZNh1zsSb5RuocK+gjPr/8Pf8+QAPd
sCXQqKCClNHxUGV8llAKUYae9sMm7E8L+iE06JCV0/PNS80z3bZBUeD0f9h6wjhY
NfoVLAtY2say3YroLjAfOCbdTnAefcpc31s8ZXPHXt/k+OhPw7m51/E2Dzaf8K++
86GtCqNjJK1I0NFpLSCV7/QfaiTWPnoHtG7THONCePzxMfitZcc8oFrcbMKCRymE
b7C9EsSEa5tSL18XcixTmfB+JVA/1+IEkJlYMgjT6n0g2bxljrCFxaHOKSA0RZib
rX7PcEDfJZAmC/YuMRMbTy/vkXC68EmV3T+Xvz1lcLosXE7HpWslWgCKT/gRqgx+
T5ZsCEnLz1ObR4qvyQFvUCWbxRbTyTwlGPrD7hYDUYNprXxi1AdFeYy2l0E4tlJZ
ZoQ3pvZ+GTvebaOrrbPPXaJMeI/zZ4yQmuGh7l2HbnHJYEFQTt1p1hTtzmWNmSP4
XK42oP8bY79hLH80d+sBH3eOCO6o0nRcoLe2W4Q0MW959SkUCVTI/u+BeirP2Juo
Xr+voehsZrBHeotzLX6IRMUCpDDfhXNmpaAdITnyNOhhrhiEAYT4vIGnS+HltiKu
Vt/ENAmJIL4HdeImjHW3641Nt9nAXMkTDmY1Ygb3gTj+LotEXAeiR9qeonrg+o1q
O61+H+jDpT9aQ46zFxwHMCXYdalQjbuj7kbIMViSdaEAu6qDhvNumPmQkwdu5E0A
SUfwrPNIl98v8B83uioNhtRmCfjGvUjaLkQGZAwaBM0dQtGYzZPftxfvaQjSERWg
6Sgq3FrlTX/gWsg5V5CIhhlHT2cf108XkFKBssuHMnSNkV8cGJt/Jfq65ah0xq5b
TmyMinfLL9vkQ0+MjadnFsB2zhchVSgc77cRmOg1rIhSwRdGB2x3vMQOCsmAIXsQ
Ti030NPGl2UYReh6Sjffx/7o+/wBOs8ZC86dmaaF56v28vOHf62TyGNQh3SjThB/
TX6QHLFtQMXu0CRo8YzFH6Lx5KsUbwA6BQcEq722z+OKRbBw2tj6d7SHqhiIPoN8
k7Le4lZNMP0R6Qy+2R+iiHdCgEN+Hy5tbY3ui4BJo4BeHs4wyLkQ4ZzHF+m9zGZX
3/uwSD+2q+UFfto6YbNyPzGMyrFddFEUVsvja6GkPS/kyvgTCGe3f917Rr+UsbgW
BUuFtYVhYRTDx92kkSdgswcEzBmngmgDGVGt+iWShNyGM5Ba+OyqgyN2IUQ8mK0d
NCVJZ0xQg+XGtFYjZ5OESYRTqFDG1EZMQUcGCrgWKbR0SnNwGwKzsbDbag9IWp5s
bqn08D76nYt7k6aT5wLlKnwR4+YH4rwrPxPYfyEvik9cUkGbpLfwEKkV6kPa7hMH
viDbGShK2/wGDbgnvSBnA5AGzMHlRclORHx2UN1Fi45aezOvmZopEmUykaauV8p8
f0cCPzRq/D86fK/qa7n/zRofSScxwPUQpC4KkpfUXERqkPXqYvftLKkSA7uvJJSP
H3DZ74lPDBkPiQfFREnjcQEenntmcbsKl26nKthBwYN90XIsoMo7xGm3BnlTZelo
I+V4gK7CYXK5XQX2v1WSxx/AivGi2kB3C2LGK26vxQLlEhak1M9vB07qqwgULlBU
d0OxrKSb7avhst+3KSuCHgxUHa9nX8JNPaMmoklXN/+LjgLhVgaSH2PaQlPXL4tA
bO+pydc806ZaAeTh7OgRcHY8lLgxI3dkfTY+8vC00EyW0SZ7QiLJnNZlM7ecj7Lt
NlVQ/8W23G6vZc5VTM1V+Y6bjbMkY628t/iXu8Pl+w/5faMRYpcnvI3ezrxYMAKn
SWcBqnyxSKLpn/XN5kmfW1H0TiTH8CO51sfyGigsiOCTMLf/qZSYF5K7fOrkfPAn
qmwCUXb2gFpfvJlacC30dJ0C1pcORWyGXnRbR+P8DloIbN56UxN4xcjLFbB73OT2
QNhBy0Vz1RYMv0bZEi5HSeRfMf+okYqOJvUJe4TOuNUdVGiyRkqt8STJyXS8ACmw
DVt2v0YqnT0yM6MwHG5uxuKgFXqaes4CPobC63yea3o9RwZ5i6vwtWBx2OzGzchG
dGvxRT+r9XOmAC46lDW7FeEwySMWTA6YSiApa9aFCJRJa2M8WV3vjE5gr6nMUT0+
kg6Nd569vf8wNRK9JXUEiHGis30hqO19KV2LlZbli9ntGFxchDApC5u1QclopUXi
MLqznonmeGAC4VM3Ck3M3DXJScM4WbCYvMMsgUcDqmXuxyl3oHQkmla93EIPEq/g
rHjK8GXCoeFTjGttRXRB7RIaV/gnOKPJ0BdQCwuyv4B6EavPua4O87mczj55IG81
P9YunJylwZZdKZyFxMhhiaK1BMECKpOnCdE5AM6tY0qgi5esQOJUtVdz6QvaUHWj
QkwZCXv/2Vgaq7U43YznD0ju35R+TGhLTZKzBW3m4vK6eUY2Lnp9An0P+M4ahyoh
AJxNnd6chgVNIKM2ZCjn9QxtbNRK+LThyR5/gSWL60W3WABbbtSO4qSZjD+YdZ4X
2iOjSCOVJ3R3+fXRN6vi10rro7EyWHgUNXe+dyMB167zvSkdlaNHlm4sEPaOxY/8
v/kgQKWwl3mIJ2JWOtaQMb5tgAHcq2XPbHd8X8p0z2QOZ+RokeGS2B8cK2Li1wQI
Syg5cf/Ybv9RVLEP1dvu+WUmNvVZCzJMSdp/IakgGjzyT4HX5C5NwY1vudNZ/gdE
gqCjb2N2MeTMjrZ0T6guXXJOOv2M4sEFGP1N0wJked/cjEJv7QuAc4Ar1eF07Ja7
GW+/pNi5+20e1omum4tABBWm/hGke9n4LcncTX1FkM0cochU8Ug4TiD6oF1rUjrH
z2uNjOX1Obbn64wKfQ2WM1oQy7D5w90vfAJ0f1tlKmLUqBuzrSs1wqkPi9QkTchH
iiO5dbwDEKHgb9zGRASClrQnzOygEGVUuOE9HACP1ZBxP4t4b9DJg44WNq52z2UJ
xgsp62L+60dD6RS5U7HjCOPQnh6ozo+nsODbYDSTDMeEj19Z/5oNPPYZTJHXFS7Y
qgF0NhDPoMae51YIRjyU3KQ/cOtxRE5wT5uOvI87ObiUslOgZVppITQYqGQNV6/1
v0XKLjTZF+Gg6Z70ir29U/DuGyqyLW9OJ/X4hBoXVc/GU7HjxrkB2lPZsrZkSJbW
++l2S7Yl8FKiMh/lxRW1zQwYKIM/9ODVQLKFRGE0mvWM9L1aoLfap8MWal6ziBNq
MMqGBb//dwvfGkkWYIK1PC5hZDlNz09hdCV6eLxps9lDzjG7m7nNqXTKGbQ3tvV1
bJTywDXTvbwnRWeuDFUfCi8KizdQY7zwP1dFC1ryBC9aLRk61pl4BkzOI42fTBLv
vDLPwh8AcdcbCqgZ7ofLguj6KA9Z8rx2zyZPY0n6637RI/yLObMzn6UhcZrU8A3Z
hvJfJgh6k/u+9ilSw3Tk0uYD5B3kzBhwm1K++8SvY4HjbwBpLoTW4z93s7VyX5Ph
D5jnciZ87Glt2kagCgzu7/C6jZb7zWqMZ1qHEmQDYJwur9lgkl7FBBFSAwx+Qt3f
rLqz80eFrJK9rjVtwVX59dvzXyPaIcVGjK0yeqVC3WgCLutT4s9FL025Zz5IzfDW
mWXRVK2z3ZWxr6W4CpxGfJgQPGP8J5JaqkK/d+lNVcO4kB4q1z8m77vKaH1699t/
8sqbw2KKHhU4cVmS+Mw7o4YdzZBHpCKniMoJm3vrlb0NKowIPT1ZPkvMsQMEJCX+
mgMDGPPx3YDrxn7Uy3I9/TB+64kvgF7ym4uZBSoctnd9/SSe4EYznCCIQ0X+cK6K
RRjFsvCEdsjNJ5ZLXKdupYDNSedlLM0TczNZI3SI8eORUmFKA97gx7AJB/B9kytG
Stb7Y49zCwVklUPvp2DNbqHPQhBmWeghSAGAUTNfIZg=
`protect END_PROTECTED
