`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehQ2UldmTPzGZ/iuc8KngccOxfiZmhxp993GEAbUiYvwVggjy8v4gUqxmQnN6N7w
jB62OihznQo1Tn9+pz5aXhQk9evjTcCYVZQrSd9FV+on+lOer0stZLHZK34S18wv
AZn1to9dlVPqOTcP90C1eOIdFevFz/6TCdqFXwrJJntoG31Y8meb9kVPAmS1TGuS
s4B1WaI4FsCt/U4CL3H8qSxDlFsUm8dV+9R7npIFeq9lx+xBneaBdojdPUySCkir
aHyNAR/po3Y3VromDzrU4c8r4ce/C1cLhvuPAHKj7EFzrHzD/jMg6tcmIOpk+GM0
FTHhkb9r9vAOMYAUT/UoiN1hCOphkf+wcvZsEilstnzwto9mAcC8TLUmJA5nH3w3
21Zej0gk1DrA9JWnEiotuZfLjFHp61ednSyJD9i4YGNScF0Ulf3DjkySHSVknyoO
Q/PXGYevvI31kfD9Qoaz0cshFHol+lZct0hE8t53Kbz1a9x4uoXx/K/eLkyFdk2C
5PhUAa5Vv2/OCOL8MYOC/ylwobtj+HMeOwjuE9mWOK1JTZl+06QlBUhdbbAuog9j
9Za/K7dgl0/As0JhLAzPfX9jGZ5YvTdeA9/EDSgP+tFRlaPmokqJc6qZfO7SdOrR
MQLPbLsP2GJLzyRP0zcm86Mh1Xw/d5AZ3k5Y0YwdUaRe6v76Qq+LdbMo5+B+gzlu
Qe6YVY9edTAYL9cmtOswGa7V3cdTyKJJXARMVKmuqKH7+9PVvMuexYqKHYj20FZp
dyd6fVjxnCvNEiz/Dk+plGTL37mBVMET6zAD9nL8ibrqkPOxw/E0+DuQ/SnKOTWo
TsxKryPp3r6m4/4TE0P8f/0MU9kMUnhZvKPHCgzov/N65+LJqTJz/VtgtwubxQUF
01rHLw6wRQ2bncgqsqgG1Hqx5nkqIoS3RmD1znDrPcQeXQ2gl3+6dHcFVufV9urV
2tb2Y2O6cduqeue1FyUMceHfDaOnb/fbTfbl7LTWoUDyOp+2NVNtG0hldW94MHwl
XLv8BJbnn2lg2zr8XUZ3SY/c+KKOQs87bXt8CH/rhaEnU0yewMvgPto0hVH+MAzo
ZW3oV+k3RW5un2aa6kMclgOTffJiwzn6nGoJ+v1UVT2CzFGknKJQxT2mKIouCk/D
JtQdpH0NH5n4XQRb+8Jp5jLM03zcJQgUN8+Nd7t8fsLXJilCWk/isWXvh6TOf4Ab
sgZaj2fqgKbHUGXlhsCE+rwjlj8Euk9kObFLkJB6upQSYqLn39CY3hZFv9J5rV6H
FINeoGwfjW3SnLwetEYeo4TJLqIyNWqvAB3lylRgCKldM1fKG0gMfEIQUWdqZiFx
P3I6AzxkCQ65KoMK4KCbOBobypq+/MCvy0/Az7kxKkyBvOiz+5aO6fHrjgaio0HA
FKBE/AjoLkk8J14FmVHEYy8pEzcGBaRfepe2kK6FWaRT9gKvWUuyd0c6+RjBESG3
rlwQvrvpEQpz7/PiLmB5NoGljNCeZ61nzi06uaKwYq8ltsoK9sunF76gS7bnt/9j
Dv70C49Liahmp9c6b3Bn6kKYyao4isu0vVuLwWuohNJJIKa9JAfRt7+vlLqLzKP2
7mG+Z+3NtFBizjinQgYgff3GbgclZ/t/a1MHD0UAcxd7v+HbJPj/zlzNcYpx8qe/
EOdW/yT4Nmas14CWwvQ8idSyFRcAIsfjFlR0uyLXT4k1hS11Rlr8MliUMYVYfhnG
GJ/C3Cz/o6hNzl0glIDYSnHNAKgFtKfhOciWuOo+SmcMFcJkIreQN/s1rB+Zv3j4
0TsAPUGUDbsQ6/c3trJORTetUk9ujtVa5YVSzygrW7zOYft+wb/LlynNmFaPTv9n
mLw7SdU4yntUej8ZNDToy5OTxG4x+X4iGKEreY9bvmsuH53LGch7+9hHCk1hVOJb
1tnNNCRmagxDeImrhANoTpNFyoPeWqJXQW/iFGKihT1G5Iffkhta1t9Hree0SrQl
fWzPH1eyhg6NwxY+ZSCEr97c3ra9LScSG0HKT3RdF2yoF+lylMPN2WWyTi8zFFvO
ZTBhGGMjt5GXFyg2CO6u/CZPRZy4eeaLZTcUO9n66ceFvH0vJmQV3vPutcs85SFY
Cd3kRQ1Aes2l/JJTk23YSMxOcsaMdz61hmm9hgz7GhTAI7uk8ehZkFWjEnfIyZmz
i12Yi+iwh6Xw/x9f/ch4baC1Cephr9ysJ5rToOfEUDJOHedI/SHIlczh8y7fG8Jp
shPWGwmCa2wpmRx8Ns82yg3MRG/raWFau6jsr0I08V4vW8ILoDzTbsRMz9Qf+rfX
fzUohmBlhnmm17UK5wUK0rxqLILvy5CaeCvuvvJtnmaLke6im+3JsPyHvl/drgKh
JFAm6cCUmdX1lkQBfkz2LU4MTu9U2ZotGVT2D6nymlMfTs9XYtsWgiWBVwXR1i54
1dkSJr/buKJ1hyJ9Ujwo/Zf/oCikhfZRZL9NqdYcnNb8+av3KaQitN7YV6KQ+9h4
bsK8S+Lk27dNpFCEEgnK9XXxPkR0+RKqR2n2K7JZtarOuVH0/MFvlsZojAW0IDU+
TkyM0rLMjbvDRwpT9KEhQNivoDX1xWgfClxNUY+8UHHV5W7yvslq/MLnQOBZF0MP
3mN4KHo3A8Zp9UP8TcWWEf/MpwRKRjmYr2uVGia74CR1C2/WCmBNoAuK7HTXj/vF
pZdTZmH9Jdx9r0IIspGoEoJEJW2jwwKZ40kaSxb0MS+nfqAwZhJFPLxV/K2yE1q/
Xb5xqPSVtTBQUHfGoQVnACxqjAqLK+csRrF6uNbbibkqmQBHUja1yvt2AuJIhu41
P+v04nom8Jf2tUJ2qcCycAcOAPfAI/sQuvulYsT7j88d4IGncRXWXjXgjzvEdtMa
iEeZgcUZveVaIYsHssvxDAwc47eFF/Rc+/YIUz+HVm8NRrNdolsUWM5qsFlsiqKU
ainTJMD3Sj2CxNMNUoya6CcFLvalNNCiN5eIi3IsOBdm3cyJCQDZZS9hAXuk0pw7
Csl/yKc4105G5RI9eeRyftR0H7V/GIdPuLYzo8LrFZmt6KZQqWIxrmHPda3QEmxF
HP9+tQnvma0cMgET60HACpRA861ay+HvaezdHxfZE94B8dssTOKzboOeJdFjo3Al
UO2d0eTLYOY3crV4B0RZAKtyQ29sEpA/xDWg4cMzX1Y5xoYypH99CbmE4ki70r8C
rhDZMspvONnzQMdLnke8HOXFR662bTqwcHLztZi6xRhzrN1sOdvahCc+lOM8M1KV
/ywibEiQ/NMRpOeGBoKIW2/bsNUcSrgrhIl1CHxAnGDioh1MkeQ52V4Fmq7hWt/l
keOB3qnLt1YM2/Vp58pFmPAT61PI4UjkdNPRea7UEm3jqwehqTl1NOso8sHzMZfu
2jt6sdZXMf4bvYHwIXWcwie64N9hGN+AczRqwHY3OY+MHrAXwBrmNy7mBZeZ4+1U
bM/I7VOz+jbJNE2OlIofAaoOjJdrZG5jJYn4sN6hrJinJly3SmRFDoLRYchs+0Pe
TRWz507h8iBgHFWo9W/vLJKt9JPe3m8PEpPoXdgET8/DCw2nJg6GRxjY1u2Ii01q
GrUDjqHlh8NJlM2yI0A/YlVZpFkiwFrgueFhpbniwIc/hlJMMjBr0yMmLRLvYdrD
9KE3QV/jQKGYnUYQbwWQ4zUzkvG692DxDSuc6/l3/70bS4Sa1EkbHSq3p9N6WBN0
LEtPl0DSPVFa2bLtdrsd93N3p0TpxAzE7W+ybmXUkX8ttnIa2HQHEiq/bvKiVutA
qgKJP5lpEFAYJi1VACyBrupamysUqFcWm1X53YzxRhK96gBUDBT+KBIet+QRidNp
pEMNrwToirXWOOS0ffs5i7CWOcHgaBHDD3F5i6/dMeO0tq3n20m+r2Qr2FO3Q6eg
Z26glZToBKiCcWWna+KLaO1MZmnC/p3lQ4dlB33Fv8hpkAQQq6W71n7hobjSj+Sh
BxAbBg9HPUvP1545B+FMuqa+Id+u41HF90JncxLjlMciEk4/abYv3mKIJmoOVFXz
1fMcbndICGnrdXt3oGOTWsi1PWj8j0v4Z7yFAzNb1hUWkn0uUVKgnR2BCY/Px5mj
JmQ/eXwwciUZLMnr6K9E1yL/S2yJi/j+qkJ28uoiia2ln7JASuuqSs0xCraVlP7O
uZI997CtQjlDSQSedEICJgGym9Tx45vQ60xV5MLTrGt3WhyuhmWyi5zdwTbRS7vw
enkD+EfzU0utTkTMHRdeXtLE47uzFdNMYjJojkfZx/UkrA6iQ2Xdj9B/yfzaoQnr
jQCaBcs2SjICL+M5fraUPbPvlj0qKctrpu7GnaMSH8iycLUNzUSnheyGuhj4Ua19
zRmvw8fQFzVnhWuumYgzL2KXCzUSTuDuf65yIwQyY1psT/uNm8ajLjr22PI4guRa
O2MbY3Pyw5xf/aH/rBX+FXAKEnlQ9QpKbqZxk/agZuIeeBdy1nw6opEJCW0qkbI0
Qg/LDy9Nf8TwCsSkZuef9dCx+sh+ufp/C5rjA4H1jbYAJxCN/4EhGwPmEdtZLXB7
6bcOXfhEiHTBgWETfPwkgWN5vJt5ABShF38cceejVoWm5znFsnqOfTE/pjWpKmNH
+WFyqx/xtyI54BrbjxgvmXnuCrHGPwToMsr3Cs2/V80X/8/QEtM/+aid1i4e0B9D
gFq+w6dtNs66YJWQ7Cllma3g2y7ykZXhDiHPCmWhJauQz90eW6cAk1vOKEj9t4+8
E7No303z65ws5zD5SiDLvT6j/bCAL661JiuEAz9YF2wLQfRjHHYzjjW0MZaq3z6T
iqC3XQdXGwPKvcWJMcSmAqq0P9dCzKiGaWl7CWPBeD5RpBDTv8T1m9rIC0zeiIpJ
nWeBNNHiYWS87WHVi5HOpjNekdi05CkA8aGNgYYk1CXD25uzWW3ErHLsTh3YHNon
oGLi+ExUF8S0vE5f/0m7wk+fFIjhzY4xxmW+svBKupE2L8xsiWgCuI8+lcgAIkyh
5Mu0DAAlDYuj9wfjnbk0G55R1CVk5VN3/OQijPe23eHXS6K8C52roNoC2G/r4bjG
SPpLNsV3jnlgx0dRjOCQa5o6GV74zuvr2wqkOvC9P3Fx5FzC8sSuRt4SVO1QZdxu
fCzwkCD1hjl6xl8LncXSKL/Y9zpHBGseb7P+0mJXCGG2nqa2S3SjZ07AVjz8lo7O
kEG1VVcMtO5mrkh5ma03i0goAM3Rp79plvHQYSmR/leqNIBhfAJzMFbUFrSXYyGZ
/PKNpep9qyFv9LVCmogr9E4yH1yhHF6NAiKMwqyTj+RZh5jn8QK9VbhVJ+lqesrx
RLz0KWoYaRA/gBN2ETxBH2JfkWShpmo8XetQICWCHe8QEw5ikwuUhBcEaJI8vv6j
Uc+EgJQEmc7RAwqde0nKdQiynVkJHI0NWdeT7yRQcMzEIHyL4QlJIO9oyyIiec3h
VXNxPs+yfwbFhlFWGqiG7737pnPq/jgdfjMonC8XOoh8liJx5wuaIaEYO86k9UWh
s5XNEkW2ZNe9B7fkqt2lbpllkU0xCO0nc1shuUnrHMDMa5W/SJUWaUTmNSM9bndh
OMCgSEgyEX5fFcRO6eKF/QacCA7GOMN1D31HLQp4YsDQNWLfmizDiVZbYGHQK0n2
OTKr6W4SgdLV+bGp7LbkAWu7wXcMN5ODnnkTaPGPIX3IpQr5X4jLCePVzwx6QaGD
KCls2B7IOZ+CHxEJqkikPxuMIrcNxrtxtjnYPCp3RSBF6AZjlR02v4GD6cOTafFq
1+RPS6OOxBkz5SbRbGHNxclruLjqIJvGVJn02NZUGMw/cuXt1iTddj2yP3GNgwIz
L5C8+GmcUBUWSAmTdYENBAzT6AmvINqrb4L5MOr+7Ur+amge4oclmo9O3J8BfWKA
iDWt2xoLuaqfoPBX0JkP8YJG5Tn6HneKcf1R0bGrSOBKHCxoQmyqBRYvQRAKTkpY
ykl6pcA0lyB0BgRtdG6NReh1C2jAdT3uQ8YUXE2FRKjR9WLPW/9QBT/QbPewbQDe
veL7X0mgbiZ93Y5h1lGPvHGFTRAZc8mXRVx+WEKjlzowcXOKKCLEo+57Z8u0lvWx
+ZAkO21ZFfLB6TBpaz/CrqkjDPb8AvGBt37JGvira93O5RkxD5wcNe0ohHKKV5Ol
8hrF+9x5u+1U5keOBSX8n2RiqwuQ+ylKy29eUwQ6SjOEJ5XNwd2il17TwzpVBk/f
3KWeUu27FKnXX5vNXpMBm563LozuDipb8Y88cgnidibX2XSKU/LeSTUsY7vy5Vzj
g+CttZM5ppafBoKDKeEwm7MLhUQRVLechqGObrD+3LeQri56dni06xMF2XMp1Ehf
eSAhLYZViDWayQq73fSZctxbORnePftdr94JTtgrVcCZWpChihl6/w9qb0WEd6LG
iIEQ1q1BGHuBzVDfCSr+uNeYJfMrGs4sfRBnOtaOt24gHDFGIjibtJPe1aa/HWcI
dGNyyNOKx9tK57+XCkeF/HBpi7eyDyDlceaEKhlfjhUpdjhIclGOEkeV5b4Ux/sH
ip166nc/k6sMm048F5ks6+u9WUlmmlhdYxEEYpRWT/dedMl4pqhbb8TYN91JcWQZ
OG/L/FdqMP5iDt4Ja3+bhtioMTqzLYNyt3nA1Q6rWkKazm8d9C9B44nWyHnFXM7m
Bo64ODj/sEF82sATHE5d9P2YiMS0D0xqn+/qAGChcieH+lgu4EBn1YpUdsqcC9U3
g42DbnO6jGL1gD4lz/ntrnbPU9eaZ05PKBm6BBa7ApkP17Z4a8LikwqaV7z5PaG2
6ecNZHGfUM4PifW894uxgDmOIUUhw+W/fpcs/RWR4t8AuWUYDwuJHuL1DLdp6IFJ
ENS0WxXREyggMKpAkuFQJoTXlgL9hpQ8CbjKU8C8QfdJcTfBW5hs9u4bZbBZqS5t
J4t5CubVn9EK5yMuDXXUaFDQ0WVzAFBUtispM0jBZeBOzW76W0ENLRZzYhkmkYHe
6PpPA2upZZoTG50WmZ8yLl9nf7gxPZFZP97it9vSmrb0BkfKbsvclij3FzySaxgd
7Dz+lffCs4CI9OKhYEi5RGfGFNJD2g3abETqI94uApsIpyPORgy0vL+CF8w1YvIT
EUvnwh3SuKtWSVFliKgfdVq5tr8jvvG7fwvrW8e0M3o2MYFGCCDssANkqyYdzPy2
0PA+WTDWTjuiTlLeciEMKow93smE/rEOCHPzdpNlDDuwe5bDdmOZ6AmdowhjPwUm
iRxnUukdQgVL+81SHGpKrmfKfrsSauMLJ4kaci1D5Lr0JqG1B54VpbYPc5/OPrpW
2lFhGWugwv1JcfHSkt4ryYL7w3YQGYUHlJeIBSMwDawupDGk5OHbo170qotrAyGG
VtvEpN+MZ95lwdZQsk9kKnIEhibiamkWrCp7qjAqfVTPnlNZrVhpVY+9zhA2lWde
LnLRMUvpxVJQrrw4Ih9x2f0WLZ5E1to/afyTKPzYd7th7PiLVMrqq5bZ2AScEyi5
s7Xm5M8ANRSeC6veVDPaACGg6VGElX7mVt6fjYz1nzu/BmuSkEVHUA4611pHxFOr
G5doxp9vGWTbuhllr3pSV2LBqiMzh2+1tL5Weyy/gWrtjvrNq8DKxmGo6jCn/U03
Tp5crxsOJwWD3zXWd/EimAgZ0o1U4VwA6diSUD71eBIgA0OyuyNtVeWv4VWN7aJr
`protect END_PROTECTED
