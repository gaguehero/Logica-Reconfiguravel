`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uwEXTkdTGemF5YJCe8x7mQrWO/c4g5CrTIyajMrtfdl07TphXs3pysPMuiIOvRKM
ltuFV7jj+vYe1A8wCAXNgHh9Hzjbh30UG43ltML+jnUgjK/lBFaSOr69mL58UE8p
MO7Jz3wpcM7nJVbkw070Zdb2O33mqwcEGro7K5K+o0gX8fnjoyfPUaXf05+aMepM
6iV2qUWc0/fEitOVK5Nb7gLG6pI7yV3d0frJ/yTDno8PKzZDTqsfTkswYSfzARSH
dx5dmTgxUAsEMuUGs0n0Dk0H+XUbngSHWvPHldzLCL60H+HVi4k21MH5tdZ/ONxc
dkWVG2Jq7DjuJO3TRJeECWVUU6V43o9gmrM7ZnibAs7fI/JcH+cic/SWgsU8+/p/
1Au8YeECOGdPTxJiJHHqnE8IURS3iObrXTNSEupBaDWlERmEc4jNOKJEAo3p7a/m
RBz6ZuMULX/zM0UMo8KvPpe+somjgVKbHF0/6j1Z43hFs6P3oErmkwzAl7TpGuR6
EHX01/5QpzAXL/GnIx9u1Zt6bq4XBpCqxI6ZJ2oHFq+dhfJiA2aEOJFCgz1aKqqY
uSQGLRYQDbyiUwmaz6Z2noUkizoGPifJkvifndTbThDVfC4uOT5mvQGw8eC3hqE2
mgaG+lKaOu+mGneL1QVSySJkfLsePZhA7l3BYzWff+Qc+9OIqmNvtfv1YpkgewEA
HllRnFFXP14wE1BYG/XLbaahG+2nnFCOQPXm34qRXC+FjCpjiqgHkTHxrcvDcwJ0
pCrtuUBUikxLBRiWUIcXR2vWi2Ere30oh4evwBDBwSu1j+Q5gBE0gdNxCMFZL/lW
85PrAD0biIt6CLWVmn47lFrOKHpn5alWJ0EBiBaOkqKaQ/wmGq65+Oby7rT/Hbk6
f9mbLfN5ydIU8qhAFYay3jgXEC8W+d2kOtPNcE5fIMkD4y0zdqMagwoQgoY/7hVi
BFCsTKzENONquEmQ8VQIUpLOcA9PfHk8sh7dX3tJxbUQyxK/oeWtfv5Tudut+LQN
89no5jmI2b0rXsjSH1Vt8UWHBEEF+Fmnq3mWpqkpRz6WPlf0Mmi0bQp13lOUQH1Q
m+GGpEgTGMBOKOxUbzff/uslIdipHQnL3QFs2ajK+RGF0cRxYZ0qJD4rw3wnPxG/
1SLopXQvXmnEcfuM3hh8EeXjdAloIVZsRWVH78LpX2tfSV3acyJvGLWhuMo5BYNH
PX/AWj1HwgI46c5Jp6DSoTJtpHMBMkIgebYmIgnD2VF0yxMY+WxB51YpDL9ZYAFA
FrHna2rocX7YHUlU2ORONXu2MdSvPImZuFQrni9pnlbz9pbsTAt6m15ZKHnnIj20
j2GEdRIeQ26WlpM13oR074jDYjVvEdRoXIAiDRCnknEbRhP2RV+Zilc9jO1CEXkz
rPqsw2i56WP8qFZWX/OoKyUW0p4eDLIS2EgAnjZq+3xjqSjAhGmoNp9VNMlXqxdR
PH+7JVwRIyrLPw37u8CXUUezXl/2WMUj8eQ//I7za7Ktnqg8ft6g/lwM+JjtTRTA
GVN16qikSSdx2bHFcnngg/r4nKxHBAepHKjkRKYoI9JZloeUtbOVNxgoH1eGvTlM
KtP/U5eWzR7iTyneBRSgMH58oIOq8XFiLoa/wKv8LZZrt/c6lIAE9HNJnkXjxCP3
mXVCvm3eB6UKgMvBbFDheGezsCbREwfv9U1f7bjr4Urlzw+xxB4+C5KFOD3mPwf8
4vcwmu+5ptY1VGLU/W2E3BvDmvF/bHWRs4+N4023xrQ/8aXBL5h4EIxvp1XBitCq
GrRyyohX8U1GdB7ilrrRZxdGc2ra5d6vqXPftf+p6oViJ8kxl6deKZsMmXQXPjhm
cXhVpDJjrmUcNNO4UGmaUh/O8q3sKLNPgygCc4xOwHArJKv55b+cZBLXuZQbQxlQ
9wgcg+pn7UyoMW4/VPq5Bj6Of/cyouNvl1IPQvYGL29Nff8c19QG5XUWMhZT1lQJ
k2eWxUNafRjwEZBDriyZHcJdkwjoOEzcDMIcWbejF0BCwsQzbpdlEkDcaGxhHN0J
TVzEBiALt9JS3MnRBuLQcBqUUHbaZUAjqctiyt+9CJBF/K+4NQ+RSfcBnD9+tHKh
C+XHBJ3svkfccpo6HyG54BGHhQxHx8nxXOikXUyF0H4Ffc7uA3g81JxsJ9z8Tk9A
ZXoF+gVJHbiCVppkEyAAULcVAjKQQZZ+MeaL1xCnwgKDBGiLYqj363taPAMM3sqO
Jx7x8lnDl0u690Fe/SHkWQ==
`protect END_PROTECTED
