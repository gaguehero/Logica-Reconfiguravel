`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfIOMDzO1Eid8WuYLC0FNUTIQKuW2VHrfnRw4zQK9KVnEPMr4GF2LHOc7Q+6gU7b
PdPD8Z+baUXI0YDEsR7pG1YxrjML+99FRyZP/J7Jh4ksgmYngMjF6oZrmO1YpVkJ
S9TsHk2AfYsCbdqnX+a4SoaExFTOXuWazynw6qquExmiQ/s+U1L8Y6MvpjeJruS2
mwv1KCmyD1zqXEUWgmR6ig/s0YQHEBmh2i/Q+vhxzbfORDggY9KBXujHWV9BDTEJ
xiWCZm5WV/EeQBXC9i+x/yDMjIJQYFCkuZwwkOZGI3NNgmpS/QHw10cCRskCHtQK
D9NWXTWXiNG+Yl7SjtwyW2BLckMyQ+QwLaDoc2MT7p3dvWHlWiQ+9R5sLDibH5DG
TmKyEwuCMrvrWbwmw+k+hhbaN3+Wjhofu4yWd2ivlmxvfj2Hgh/4CP+3QjclzTNg
u08USh+lVWwx/aRhz8W57QlKJo5Tg8a/6MC/L/tZ1aQ0vU6QqFkfRPdm84RNnqSo
RUoJulFokYJHPKirNrNGUJQkmINTTiFXTETkQJnp0BNt/KSlAv5Cx710Dihg1kwr
HLN5/sOYddVNz4E2/Qlg6rgfDH7F2rzCy8/D+BRzpTcAkqSJq3Ee/9OKVszl8UE2
a3XoGk9uMgEp5OjibMKUr54ALm+zsOpSbSfgM8etiZrLQIPz4lz3zsG1ZoafiQ/H
VXzWVfrhGOz0/r+bxMQabzwG5ctNfd3trPGgJW1NmIkqzd44ezrF2XJiHj82o3mH
BUgxVOVq/ckVKin/PwwbxQE8e93VzQRfnRltW1g0NHEtCYe+apA4mE7ARikCN90B
uOVy6wZlF/B77Yv8m5ubAi6dUhySvZTNlTUx1U6YASGYr1gYd0vpk6u0eafzGOPV
qVm/poR35ZYPGPyXVZaxOga3MNB6PQsc65QeQ5nCEWNPMgHmgzh78/KCOt9Wyxag
8R4a8FL3h0ZkoLnBnj72dslLTugv7T1lMoO7D7TxUgzXxpICPpDKQoN79CHeHtBL
HKJKmeYGd3PjvV3B5ZPkpZgHxVNxaXWD3uOe+pEJrwwrUcGCs16nq2GBR5Vx5jag
c0MQJCFFJnRRTvzeUV8DZvkfm32f4vpdABERse5C4oop74C84kCxJxZty4x7U8c3
b+XQ5ojEGCCkvftDNN0ASsYb84VtgcREp2nwfekGlS47HyKmnWnXOJBeK7fYfe9g
Uspg41hEyh6PVbAaOvA3f/tEk9gKuqaJgtRIUhF9VDPZY4jYjzAo0/cM+YfNCMrd
tnSAp/hpPxPI+TAWXeVI1buvs9erzOO3rmKKqi7YO8epT4960tPhYM/tt29AX2+1
9UJdjGV/XqJFSWVVqx0MNkPrA1T3soeylyVtFduAm9OEBbRjD02y0MSU/48FNiP/
U2SUXa/x8rJT+AwO9/rjIvWri9DOMmMs/YZnXWgBCUDZi/Q3S424aZMspb7CxJMZ
Qo/ZT7SXpiLwF15iwhaZ//ekYg22f4bTEayQYIVK9IOgnn5HEiMB9qv6nIgd8GQm
ZTtkTz7YeLH8PBTpj/2NgMQcRbaKWr1z7x9a68HEa7MX72haie5UDo0WAFhz/54n
SF9l4/CuBZHBTGEqzVzJyznAS4J3wrC5vTPnLoQn2dij93XoG2SS5Wes3j5w7wRt
joXoBHHxMO9V/SrBRVkP5wEyqQFr3we11GhDhoPzlfjPTxvBTfcs25+G/m/Vvw7X
jedxl/o9AdY60Vn6H/4RXewZcmKgS3KZYAywpRNNFbSu+fWLpY8zgnw28nP9CBJG
6GpZT6Jg60gt2tuSl/ZVeDRyUouRQf6WwrAHI1D0lwXJufh/n93j6uaxBFcYIQCh
CoHwPG6kvBLkgVdybCSb7mqz0gzCfSjuleYuAKK81ozer2yQyer1q1Q7wbUoiWXV
+PiFtXKNx9+Q+vC0CJMImgBnbJxpRnkDwi7tVFytFRTLGkZv0Gzw7UfmAAtcBvsb
hujv/nanF00H2yrifQk6k6RPerM7EyXqJWKBiZAf/657ME+yhCDtbOU3a1jY6WLO
3k2KM4MocD0uIqAEedfXEUVzOWK4sJ2BTMbAbqPb2OQHGfVFKjAf0jkDBm8oH5nM
sg9DiSjegHVvUvFzHDJP3PnEnVJQfCeJ6uoi1UzhGXiFbOiR1hPyh1MfMh4TejkC
EXMRAIm8Mq5hohY38nj0RKOnquJb6O2ymqh+cAXwlOA6cSvpx/0ZyycMa6JQEogj
n8qVVXDnDNPUcNSvVPVILrARdPXDSInkXK7AjpUC5pbwfCv6j0r9cxuTyjfgMd0c
qO+4VmRmPY9rkb2NkCR+D88TH4GPiE1Jzwr+W15ubzpn53DY7zBamhMvIzFsGHeJ
WpgPS94PCbTu1Ugn5Iyk/mzFwaPSU/hgVytpbsPNJn4Ostu7OZZ8lsZewDWwsLzg
V9dwqDkyovgEYlW0WE/56V+Mfh3EcuJNz01vz5rbIy48rWIxIrBJdrTI/BNu5rhd
4Tz+1hlw3YOMPP6O+0EbhmqnCXxArbq8VQUZW7WfkU1n2mRvKEg2pSfmc8YuiZX2
FGQFepFRrcgyOx3vOx96S4B3b2QBkgag5eEdS3RLorxj5ylkCRZwL2X4WQ8e+Ol8
Axuao2iG9qZ0WXEz2w2aqsHIqpKqeMeQ6r8yW6DyEt5Bz+HfONawUyxfKYFW+YJt
AMtgpt8UHRCVBouTbKrCcAsPOtC8bvS0cvOG02GcZ9jSMqXKPMKSfNFq+/zYuIKQ
HO7eduAMzFBvG+198sJZ1+la5O1NSb944gMW1xk6gzfhd5vDfv3tjRo1VjM/5qF4
3t7Fe7irqZPWvTH4wfLO4ggotMyj6B60MWQN6jBKzsWsDvRSxAi40tRSvfl7wAc2
uNDo9Bd+dsst7Nz8tYoI35fxUqzkoVH2REY5UvjF0swbkb3EyscJHPHs3qOT62JL
Gz+ceRDOPmgzXnPshssZChEF9VjBhBYPnmTQdmmnPAntrccJ8VqHdVDEQ3OzElei
KuCb5oIM7ZI0EGlTBdgqH+nfYJ1Xgcnen3JendMkrUDdvdYHeQIjGi1oQuvEgMeH
YUEL41F/yp7CeRlgiETPaO1hnkSW/QJ4n1rg8bVXlXGKTtM57MhqYyz43M/XHKPn
GH9nZ0g+da2uzZ5rU1QmGxF/FpSNQD1RswG3JJOxK4ibsyyvUbyMdLkt9zZpjw8l
DOlfeEhWxOEraABwCem28h55uUTFQyXJvIVicrYdPHz2wMZedVm0/b9/3LKVkbaY
wMCQMy3cCMi7qVWR6+T+gIzwpeice2QWDKeWzBlXN0plCzXLcDelsOyyxdYyzn36
1GI68oTGnKjagUeeyD7tHHmwhiT9RcSjMktsG7M5+3vCv92mkhWxcdQ2b1RB3Dha
TPkFkBmCAokH9Jzy9Ao0Vi81pIQvJz6l2lzVRoZLGZfGM07phj4uXJPghctEsLuU
tMfsoOeTiUkqBUb3dNkTa79zlPPuLE5KHGhuPxO5uWq31FSsCwgtWvBXKeN4THUG
dgducN+PDjo/gTrrOtTYRG49aLRferkrQHxzwDPMrwkAFnLbYsKM6onvLOQcz/jw
BxeFy8yPmLS7Z+tTzCw9bv5/hXtqUAPq5uhXoEZEewpDBFCatBBkf5TGgQFTxF2/
zbB1ULn5bbLAa832mC784+k64mCxKks1HzyEFtJTOSw+dEViqwEJ2SYJ3lpAROVu
va3furvEKQMgXe61P2VHbPuPGwA6UiZSbwEJg+2MFyX9/ANmCvabztudyCkJxuqy
2ufCZflhGkZoHKjQzRxtap5yGxe/aZsknUJ1Xlv6cG+1ZC1is40zIFtU7je4t9jU
uYGH3RFhaApR90t+Cp9RljyyR8aLZOUbcekiAmNonZa0umzcWxBbZXn/lIzR/i1E
mV5X996rfpNCKBQOtS11fExeMTVkqw54J9eVvlqX7BtEe5QfPfjXSWPkye95zfuJ
rfV2vopO3SSJy7Cn+XIOfzVEHkFzqe7SY25m+S8rCTpjVL/WPmxfBYdxnPm0y8Ka
u94c0AyIKL7LGaZVeCtgeIP/izshg02tnFsu3NwEydlHxlaoVBM29aPX6xE2WWn2
Of2xDQ6T7YdIc6+L9Gqvn/ckFcB1mFvOi9bLWZwag6b+pd3YFhZWDSZFPWBYrPWZ
JkKK8P/koUWTT54052MadZahhwnfn+pIh9FrSV5YNhfm3u4JUoIc8ReVg3Xj5G3p
tvjSznb7r0Xqu18HMZgaOLsT4llKkw+U0UDgswFPAQVqj/MLODdbrqdf57HIzqSU
hReyTbhkDHQoPwt395dfYHXzMC+pB2tEItWOQnPumGVYrQ/FK5IJVyvVSoYUgpS6
dVAphx3tqYU2ky4SPqt12LeZyKOd0uPe1zUi4TgcfSwriXrUjA9batCbO2yo9iPk
9cskPAd8ctvcVN16IHdRfWsbGhoq/yba3px3nBMmEm0Qs+9HUcsHmnHPd9ET0QRk
5fwXJFQVwm2Rd7dRGW2EBK9YhOMdvLxQpF7vxFO2XLld8gquq4A6UVJSUlP6JSWy
pPJiawazfrT2roQo/Xpdu1up+07DRWuscxxolLNHRtvBygk9PB9IG/3UbOYG4Nql
/XzIZfSgbiLmrpyGNnwNPdmKCaHmoSG/OZZ2+8/6mFgnhIPs3hS/t+s8XJATqnIF
kYxwIDPZBA9AXXyhJ1WYLt+1qpi3V8vYcT1bwmVKFpBVrk+H+bS7e/mpX8kyvaby
7e6rIYMxa4uYPKwDy+Qt7lvhncilc1S6XoPSRdJe0N8qnhnolGhubZHtY5oyrTAd
5rhAPHH7c9nWpC72lfMHGnwZUQK+RNDO2V0BoynznHvdrI1JqCpEdXqZmHafYHDu
Pzgyejc/fp7zA8DM9cnfiTErQRvmU3fBCi1aZ7E7k03aw5Rw8VROeQzdWZvIjs9A
7gqORFONQyJDqWOh6T4CsdTqo0wRpwg3MJlGKmXWvnL6npcKoLeoss0EeUdz5NVm
bpID+i5R7AjnRZRaugqlAhwK+yBtk+Gof1RWP8y0NfQatT43/8D3NnHmZLoGzQ4r
X4Euw79zmuJt1X2ys4H89tHu9CmONCp47sEvC6fCTo0Dt7b3x18TTvOiFsHBpNDn
aK52KVTQA3xlDhnlyz/Ou2Wy+L8WyLBQOqo+jwU3wpW6EeYLwtq3soqJio5Dol4m
ObKOHUC0WtFB/JPXlxPvQl87OPBjvU8GFmrkwyuwh2ljsagBGbpCJ4hndWRIAvnC
lh9LtRX6+MPBfag2157TDYu8OyKpXqapOqA736sRo36tup8+sARcqmpkKoEz7BNU
MoZF61klgjMcglvopodRywZSElEp1HAWjwsbZpBS+JBvTAWCzh6oVkos5SG/8q5g
zuAaskAzAK6j19CTMQTTqeWvCReyQQP/pSdnYP+jOgY0osNHz74ctvPm6EZVxKe8
PVb9ARLm4de9FxV4TS9cg3Gknj2lQubM61L2hODfM3hTu879QotkWCERoCdniL4r
EhZPLaOTTDTN3ZxtapC2GQ==
`protect END_PROTECTED
