`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRxCeT3DotbwZxa4AcfLwR72HbsWIGmhNkoQcZp7aigIXG0ce2BffH8e7fmkExhX
3HmnyaEKtk7O+RqlzQwfZqPjzZjmhiLTle8yZekA26uZi4CkpFn2NScvEHDbJNb5
4tXfp+1BnfmX7OKr6wmT75OkV7fByQLOMzY0sk/sOlqE3JFcVwwkrXLECWc2CLgi
I13ttCrq0WZVKRVcVa86YAziQo33D1MoUGAH5AeELA5/kVUQJQx7v7C+HvU6ovH0
LtyjUlpe+te86yXGLUkqkwbf0XkhXjVikeZACx0Zzjm7QY9WS9SsyOyD685cnMdl
e5O1HghU3HmRLoKThPe9ONgBHp/oAG3IVZoXrFuqq9k3p1/kdmd8K8t5rzBRr7+C
wRKiA2yUhF4umwfA00IP0CAqNp/C/L3NKEFI+CHasWlMvsLCvIsG7HBsdXNd3PW4
PlWMyQLCbOZA9yKpgVFlAUYaSxtnYBthanp+pYdblNc++rHFUKwCi9/p5QvY0YDa
LRqHKs3YM82L9TNDaCP3TTU725NbXTueg7hYNRxkYVmPUs68oS/BAMmUkGNRyJ7Z
aDmGYN6cMnkffDEk7sAr3zjl9d/p/ZOci4RrqMt4nRLY0fqpSnLscVIWMLuy40li
kgCTfXUr2Ek2j9PVtYpwyOnIQwJ3D4q4IFvBL4NRFViQsTxgeCYX+6t9rNFkpmu0
BezTRyN7zq/Kx0rvyI9ba9PWU3FKgVTsc5hQ5HSN5iIdFwEsLBMvvLINMDIkN0dR
ohbuwTmSKel3wTiJoVMDyukurcTQDICYBsutseMAFBD98eyimhRAQUNOqtN2Kd5g
aXqP62QtRWQhwt5vfz7Nr77AlDv945Z8794nCiSGNyTusbql+y186i0q8fajZHBP
PaZQPE7hZrp+6SNZnw0LjciXTl9ROsfu/IE7wDMQ4vA7XevT/9H3EYTFCh4r1TXk
6/F8bmp2e/D1QbJr0SrM1akhfeu8pe7PIxV/q11vB0bioAS1HrNRObbN+vk5vGDe
ti4Nutc/luz9Ko4RpOXS0v2NI1d6e/C8x9m5YboonjjeINHHDL37KfHEr6f1QVlL
q/nLD/ZGfhhG68q70xiTlJI+ebfbfPeUWKhoy6U08nGDKMqB8BTFmWuKbjXJYlvc
PAsk1qjx77DkurbFeai0bmqlP1wCb3CwfaNB1M/dIzk8cObKvJJS+iHG7fxoQiZ+
KH1jZg5d+3mGbCF03qTW7pLkHlYbTG4m+03FRcVx2Uk=
`protect END_PROTECTED
