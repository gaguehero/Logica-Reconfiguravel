`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0J08b9muQ/G7B8Zse0TJLBDc9FutxX7HwT+QkI6sVyMHtTK554E5iFkrHYfySRj
I4dXpeVWppHNnBQ2PRV45RAJh60DktywHZdZNM//iJd/lbhoKeRaQRX9AHf+imLu
HKYvfasVa3VTIqnrm5czSflP1Q49SAX2OSIHnADSFNFouQGIWrt/nd63KHfRrk1c
No0jKpTUxN2W90zlybeWfsK4Padd5IyFw4oaXOQg2ViF5y//FCNZkO06ABA1OzOY
YBDu/dvi+xMvmecZzAKvr42rPO5NL4SN4rCQfy+e+8gec8VEkg5TdqlIaj8FvB50
hlhF85E3ZdWJHc1vVCXFZMovXmu/zTr9P+2Tcnt0xK2/ZQm6vcOIgQVhoxh4m+tN
y0rSTcXKvNfZYUrtjSOYHnMNRn2+Q2bH6K4j7e3cHPwb52LGK3CqJW5xFQSBKl1U
IAWN7G2sNIuX1qLiapnAb8B9hCSIwhTJeOo4vlRX+6xLyUJ4lZrNWo408IH0tC+I
KN7UXLRrgzXNU5uCNn/hKLfBh4ukqY4ZR7t6Y7TjNPAFtYmbC3yMyNVIgO2N9ECF
AIcFIc1+H+733AS2246ZszUGqemCTG0NqJrUl0n+FtOS5W1PXFChYQ/PsCXSZCbx
Mmk5YJjfMf8X/Z89RQUDAgcl/mhcYi0Qw7J+opTixZVVPhGFw7Rbrdh3f22/GaMR
GApUf8r6OsQ0qvRglrzpK4q/RqWg1OjfWbjWLQ2mXTCSAEtqAToxXPz2t0yAZ+7c
LkKZ0o0PTirjy7XVcOyz+GUHTO9SLhQGIWe/pgn3+YEybpLuUYW+f3iAeOC112LW
KfdSWBbO9GMr9Kx0+n+1xSwPOAkkFmjEoXgwmXN5hnWYwgAZp4+O+xyM/t4FcEBC
pGHdB9ckSGEqz1jvZpv/r20gvv7IUiMVgCqJJ267UVZBHXvIb26NlKd2OGjH5Cpl
Tt2DPboVsxugTFCP4Bb+NYhIIn52cmkckARq+OBflE1JYYoKMNkqAXDK43Kb8hZ7
MgyVClNej0Zd2HndgPIPOZYPo1KvtMpC69sPDF6pWJ8fvVUKp7CmALUTaUSjtxqO
+ICGcikwIqvqY4zk+Wh0vDxSPSNF4/+8i3f5kiEMHbDZuy8SAF+Uk51huhartss0
KDSZ/1yBsZ1J4N6S7rogaY1KknZxrzL9pyywcsVICEvUSKnmPvJ2xIprtnNy5+5l
Gun1VDG9R20luobCntrK9UjSYl14/NAT7DJD5T4e9yeBYU7EjtMU12s7rN1ZsfY8
O0xr15RUNjJIfqY+P/TmnXqQ0drEzJAWY/x6y8ojUOEw7OYd7ii8DBU/HbYgEzJl
zseKlodLawYqiBJ+rffT7DQl1eqVchGOL+fHB9Upzjgn34mAsT9M7OUdsH1LxFlE
xhWaQawm6l/SyMo5GdLVioetPvuMdoAH99nLQGfevYN2yeC01XYv4shD0JNTShWB
eFUzXJj9d+CwUo63guPsqS/NqCvOCRd2tE3/bng3hLRNYWJxtg9b9hb/AXEMniRR
PhKJra2M5bedu0yVWsIyrTKYTWz/XcGRKBXHy+i1sbUO8WPKQnABSnRK9Z3Q3K42
aCPRcutMimLTAykoCMPQArpyQWP0zpZCpTkpVfsFs3JMqzSZlhpIBj4W4EjFfsy0
0fX96uPAh6m8jBEk+w9j4tqe08Wm3iv6p6eLJVROWi3sp8GvpX9RvJtQ34b3Lzww
gPvymTl+ullDoXCojlfMgrv+XGdW9EE+4kTMgGmu4EMo2gGQEt4pzzHdRDy0EZgr
YtFYNLlTEaNVUtIOlDhPNRWsqqPooV3GwyHK7w6Tx8UhqcK38Cd13IsbnDf3wkE9
QHsyW+GYMgXHJtrZn2lzB+X+f/UEb1/3MzRVVVzWB0apgBrxtMcocV/Vvp80nxeB
BOpSGCpGZjx+q9Q6JecbBiYQcj8LEJygj4K2jaSyKRaNMZ3XzwqodggpjBOl58FA
JPsoRIUeKr8UbQRFX5jUWgPQa4v3bXAUisS17d0uSIjwGbPfUBofboHRW4q0jo6T
E/S0pLONxcYhujGaXJwa6Q==
`protect END_PROTECTED
