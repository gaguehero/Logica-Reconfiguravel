`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1eiY8+ztkvXjAHk2Dv+NpcIoGFtIp5g4lPhLfmypyFG5yw9rzJFNfi2V4GX+4b0
EG1f0m8OmiUB5zWx+exDmfhrLNv5ejt2bOTMrhWMAOfUiLfoxPAwPQCSBENYE6zx
j8k38Txp5greW9jH+oyDhULZBV1d/nFtthUKSsesqFM95Pv2pU7Rx8VS8fA9t4tt
3aJz2desf7OY+wQBDLpVLevXBwfD3boF5la7AtDrrGYUOsSvYKcSWeN5mwJ+wZo2
aQgPj00tkK83Pw+Wn7AL8218URtG38HkXc384p8HJQR3F4dj5iGI3z2mqs7xT+Ds
ysaqRRKK0qjF8M0j4+tYnx7QHLRtbrfUxnXs3I/DZT218/NZ3/l/i7Ezow9XSdkQ
Vc3Ag8fMjJBw0an2xoyuP3bBWR97pvdiUda64wo1BCGkMc9SE0b9d7uCfmFxQR0x
q+kCfVdwjTOZD9Fld1exJzCx3SHVMFt8XLlFfESQwvGJe/4QuglMfel1BxGpPZ0w
4wj+XwKtPywjSA3XTOW5uWwCu6tc1RYaNK/CBOB5MFZJCSi87INzHwM7ifMVd43e
m3yjCdIoNSQt+8S2Sk8Q4h2RnA22kAplpcnhyTfBj1BwxwraZSseKa5NWp0GvN5C
ojYoCgLYpTzXi6uaq9VgT1s/ZoADUNzvL0m+Q8KxrvXu7k6MtSJC+Dd3s/+XzV93
/rqgEadigRlo5Aw3VvmOKmvhFNnCpmLrebdTvdJWI9bdCrWWFDVBF/Ztg2TK6CPG
7L+nl859Yz2vxfIv+ABr102LTeQAqiiL0bsIfke5TyBpC/gb270v52gaaWaAs6zg
m49wl9dRf5cApSvWXCUBkHeB7kbmLYvs6RcB3TyJkYoH9UO6UDPfprwcxGxqJpvI
ljG/nJZJi6FhzcpN+EICDjDf4XjyblIsJeDfpwA2tRoPX/Ka4wutXdNt02936Lhn
LgQW9sRtjEkxOVJBc+mPUYxYVm4AzHdZTGLZXaFSlt/mZM0WVFgoWxnfTPMw92D6
yRPVGzkppxUwKBT8QC2nOHptmWwvUdLdI5wtp3sXVfB+Myjf6kGSRb8t5/GuxEft
18T8qVM+Kw1RXuU9aePsfh4M6J2LdN59Y744JkwxtiO5fOXxqPVTIboFZFVlClah
It2K7wtreqmPYgq9GZvE0wNaT7Cf2GZtLJ8lVPRrA1xhDnGal2OJg9qeeJlBHRlu
p7jMqVoa/PcdXqUQDf7MynVIRDUHNeJAy/RWdK2xx0ea1btAuXZ8X7AAYZu6DvvM
Y+VP2L53AsSoyROZH9Eq5b27mG7+pkkXDKxN+9x/CDy4p/5B+3/C/TbgrUqBV0DN
8nmjBQVjlZOBRg35nUK6TJqXQ3D2cqlbiOjzwF9FmtFDha2GT9tS5Ls6XFyw66lI
U03aOuQce9W753+XAT9IzTvA4E9oAJOkwEDxpNdJqch7fPP0jZ3MzaNStkd+HnTT
NNeFnOLxQ6kzCU1BrCPRdsCDmssopvx6HzNeMzJ4POPwgOUrr5SENsOjwVLe4oxm
5QZdFMrXFuI8krED/bUdKxLOql5wlDFz9oMXuKNi1jQM32QFzpleBfiuR1SFXpSZ
lnqotwP51yZmtBOheBeSlrg4C13rP+CY5HCnCNARUsYfv8OJWh3dh6iGR6+tQ9R5
za/Zx0s0V5WoEFIlZWorauHCxbaCsqxzuioBSdQBtKzLRt++uTYT3td3Wtkb2xPz
LqZ3CHfCnvLE3HXmA+Cb3ukT/JgQkmOqIyQQix9klryQsTC7CpsDZYEQQPEjGfN/
Mp9USzB5y+ao0/4e787x17BXmMSI5EaMVJigyYmeoU3f7B0qkIVP9Q2MS0ZnQ9DJ
dAnep9rUP2VPokDDf/b6hVC8obbopaFtxP9U98OPii7v7MF8Co98XLoiH5KR88LP
/DLElsU94yPB3ghmS+H6En1c7Xve2ycWuiK+aKqB+rwesr6jPo8bmhIaLmTb3S2k
f95Wp1HrRzjyydz9jKxpOXQIsocp8bY/9HgQOHDqvL7yT/qidu+LyaohelvUF4eu
1+ebJaz/eHCB0zdydj+wUhoFJ992mOvsu0YZNwm2auT1vGemP1n9EKuxmqR4MdLh
eS4dxWcyzO86JYcptS7jsQxxjVHheHvK3lB5CHoVEHej1wDE/c8A73t+ObBfsFrO
kEQ14p1vX1T8cpfsRqsJuaG6zXWumsGWlGV+H7dm8hY1I3v/QbUbhFcaM1gfoEYW
rR7D5SkAFZIgYEqAXaPJMzoqMOqoZS44tpNgXAKkffCibGnmHA3m7yDhMpYdEgCX
Mukc7LA/fMAZ2q18+VYfmPsrqDJwTCHrXtReKCJKTVk7GlfQhpNpqTRDeJ6RvsV1
wdy1R63J8wFpkOwHh3PpF5zE5jQ94QwNu55o8pLUI/YClfT3+HpW6+mIUK9lTbu4
7Ni0nYWyzj4m/t36fXwXFnACyrHpY/kZ8V7Pr/ILQaeVbCl0Q6NuF3L+1Mc3uMxT
W0IIvOashQOH/9eO5Ws1fp4uAXtt963GTYmzWbqShawdskeUUEggL8Sd2gkHOb4U
nI8vbUG7lGcbZCBEgcmaSBS45QeHd7YRLHnBVJDmRCeASGNYmld2hPASEsuMCadC
o5FBFGoDfEy05fe4O0Zt+sBnq6SEM/wmlSvB12lNiX1hRhOHUq3hh8Dj1jqSF0wd
rla/0AilVS6dPVmmvr9tVtSC2OUORH4ge709rvMW1f2rpKk87NcUhtj83kB8O0kX
cu9ftdd3dy+xNiQCNWm+5YoHPKvQwOEav6oqO0JKZJ8oqa1NoJjSlNYfwHjg1lrJ
O6j7Gy0mBKPakreaq5gBbQmvkWZo3zCtbVEedbl1l/nYTnZcdkopWUfsVp/kF3sk
jx0JJMsAutHA9jgzciPmvZ2l15KIMJ42GXJBwh9Bf3z3JbkhtoEI/CkrYaSAHPBJ
/BrfDeTNVgRTEuSZ7Pv1gLG0ufqLBru/hV3xc5usrCwHjtTw4gEHBZk/BOiyNTDD
TFUB15+8VTMWKjUtEFvH46Ue3ABz0X8L2/+8qIIh/CRU/0Fa+6ix/B4QnqHujKwS
6rAhbz+jCvxeqi+oh8a44WDgqcb2p45oAg3oQ24emYwRVRENKp3LjcpO0yClk1ze
5e8SBHFkGoxt5ilBwvgKE2JHt8io5AxfbAU81noaZDjsskqJdE2Y2+gRrTHuQTuQ
r6DhdUVGlAZc8hD3WPoWBUUjHMTMxGYyfrINlFz6eExTIGVowi2wni8QfPv1sr71
n5OTPf7rxB/cfje0uS6PmWSfsXPa2RQ/+jcjam+mPrdJ4hfhTtvjilDlI4lfcnTK
DwxBbiluaezHPs4wVMsbc/7W7tIvqsMEXaFIaduxV2RI8Z+iBl40dNu//jYv/Pg5
2Y2i+DAvYLBDD3685R8uRsGl7JaR/HKr2DDOoLYl3NDQbpiURmxNouBpy8yNt5ax
xGk8ihH7YQ4Udp+2SaJsmnVttzoy4PL64t+1de7ytztGkVsWvlo0Xzbte1KbFeKn
m8aIaGjTI6MRy16xzULKJCjTYYkEZ8+kUz7iYbuhgpGl8QEYK3f362bNmnB1i6QW
gX8NqhhXk4/ynSkESfyR/ZkksqI+6bVcmjOLmGKswEq6jQg3srDTUQtkz/AmlRSW
mYuSX8X6hsYCxaxMvd3nsCCzi7UqeKb/jiN++H8ouCZ1g5wZVdPZsngWJzecjryQ
KjUWALqq1NBUdkhlxJjIv+1A3vtEuxkKsgbV0epO4M1cdb/JRFpOJhhaNgTDY/ZB
SIKrmiV27jxOJ41fSP5o7kAVZIABE4N8DbRsPsJLbN8WSk5Qb2yDjXO0YbKYiAUy
inbSGBXmZqwptXuwv9lnQvBsTQqZ/6934p9vUsaduMk1mu/9ta0TbIctjkaO5Bto
NSwpvH2JzME4kEvjdkwVGyJE7rI8UImBh6Q47zPjspFiGsPIv6kK4QB1jybsBvUA
K2QXO5FZAlKTee0pH++VnQptwD9m+bm299y+YdrhwDiyEc1KBAK3wbEzX4dPfLP6
o5PRJahzUcbPNIfQ+vriY8HJ3/VRiPKEjHFd3tTOAHN8/elxhwLojskqAUw72+Yl
MhxEs07ZYu3AAYm9cdYXwAJto4d8H31gRCG2bsi/8FIR0ukKDEDEAhhg9kJaDwKH
awM+2/fE4Uw3Z4oNEwPKKYY/c0lyqm7X70L9NYWRGpjqYh9DTxQSEmail7VFV6kg
CJw9OzrEP1cx/jqHt1O1zacD5b3GBrfCOgY3OiC5EMZRq0+yEGqYleXM97lNJB9h
5B1hZnIWPH0SpcVLd472WR5mmZEIUTAjx8xXKR+/UrvukaVO3tlmBBsYecNoW3q9
7KdbiHBhT+bcD2JxuBqq2O8EyKKFjh80vX+jWHVgjKuBVGcuFZXHx5abVvK0/+51
RyuVY9hEPuUO6wwxUUwNyqQtzX+iT7iZ9pCpv+8TukkUc1E4n13Y5AvRlVSYqCmG
y03oeJN1IthT//HGLO8b4D3rUIyfXw0UAnekojFzosd+HWq57B+k5D5D12sxfLgV
7IaozMzFP22p4cdIHRhGGpvFERLcdgwO+maOnDZMeoIzJNbA8ijyaBMuD4DeBYah
dkoyYLP/fwbqlEP2hx8YSraRvr8xv/cgILFExhuv2DaXRFnAjkGVi3fUOIDiRUZI
sisebMmrKzxh2jVlOaGZmSQn0nPJAJYl6UADnuF2C3ji6fohnePQjPIIrMy1arDt
OWOccjax3R5z0RqF7RQMvnoWHXbJnNfq/HDrt5/IyZuZJ7txCFOTKmCuHyhZxslP
Yernvf0y9skq01xqDbHmA302St7JihaB45PREFd+lvmfC8tvsdjNA5+Xq/EvWAmX
US4pmo3fUNL6nWhvqYA4DuasEOPZjQXAa2l3/kS5JbUp71kFwW4QGtuoY96wmF++
+TLYIQV5YBn2/XmKobkDbSzdlMPT2NrEaU5Oo+YE4ORenzKtYYYwprvq05vdjT1s
UKVvzohyCw3zK6macM+86+kt3PfBR8KpVB01pN1kFoxHwQdkRGTufARmYL8M52lC
MPX1oY5aITFskIkGskqlZwZFLnsRFMc8QARZG102H1fdgbejmjGTB6x9dgJZj5MI
VcN53YdF+WAU9V4HR+e9IMLmr9GZAsNhPa1IMKtP78rFbM2PwHDyT4nZsPD/gvAM
qDq3H9I/aX48VWpERyc4ywY6+GckV4XLvTl9RXe64XUibj93ygCeJIojqe0OgEuy
16HGZb7Pf3xL9CCF6GJiYSeu8pNqql6N2H4EGrVi9z+VBLcEYjkfkn1JRmi4x6jT
1rC1DGcTUSl4OLR/dE7axyA3KZ8iSyZQxN43V5vwQrm24/5xRz9uR1W9m7x8OKMv
OJMnpQOXELmQK3JL19CsxmzdJsZZsuuw3eXaV9tLJjjW7edxOGLW5u/4XttNS7Sh
UnaI/9W2jG1BSxPADSUk0swtIP6gimoyOMdWpuLkQLBbddg59c+4VBXmvBAaYfbt
S17QuuCYoabnTaaYPruTRtFt0DeENVdqaffHt5qC23b04oF+9QN9Zxd22eUBqc+o
ARg11kRtBkrKePU4sJdH/JsUw4NKpOWQyBs7542ip0huPRt0ZFM2eAVFTBz9ZOkv
d4js4QByFu4qameYx1PM/dG1Gs4tK6Hc56HUFT/e80UhxDK1nbF3scmxvzQewJ5w
Rg1mLtaND+notdtaTSbu6AmH2+tkgW0cttWLymMUNyneZPTM2ufvv8Mnwi2Uwvu/
N9OLFkfWThzsktQCUOryhlBCTU3SQVZtL4dFCQPQntyazxW4ubdx5K0QiE+769hb
EypIon7N4FmdCLvzvvhdGMD/uATzXjlBSpt2l5pRGBwhj9CfuYos8GnueoySxfIb
6dZtMFcsZHMlWS4APHRZ5xBjl5ByZv6jUZjFCJNzN9Yrqbz9wzKNgDycvMexGYaQ
zy9SqEQZQy4eKHH9mtO8K8YDT8/I9AyLpgc1evSfR3zLJ2WwANU8F6aQgEThxkJX
3GyVrj6Sr1O65oXsa4BAMhNW1tMZTF0hztbGoU1tG1E=
`protect END_PROTECTED
