`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1Zdz7J3JVO5c8QTAFUa79Tup2jAXmRnM/0QcmEV0MwP1i4VbkW7303ZG1daIXcz
v1U5HaeiUNoN56uUpev70paDUQW+B0Sf8eHKoqjwWm4HM6pcz9a9tCO7Qy0K9QFM
K1J3PU5qXSBC6XHH4kUnOi4lBgNmo9eD9LWVqdRuFCDqhL2I4VDQwkJ+NoS7rapB
bXY+LZCFM9MO4kOoe8wPqT4K9te2BUd+tchK04/oGsBy8D6BVnsMPXTLD9kV8CeY
Pg9acFj8plZlm598enmqwEMQ7grguR3ZaIL/TgFe7yeeykHTdahk9EeoZHapQXh1
9/SsCMLu72egmQEPI6axe3td6wo9CHTJU3qWIj2Tm34iZEIwfwnmUSsDN/Qf7Z3A
Ox00ZAxu5yI8U+HLk1zUKeu/8H1h3PJf7WOJBAylVL3AEWkv61hb1yfJAN1uQesL
yL3x2v+mcR6s/XkllC1ErgfhFcgjag7H4up2rV/zg1kLt4uFHkBk9onGaOWoHVjE
4oGggY9C7QJRY47eM2X+nhiPMTFq1QGYgy3HuM675W8OCWZNmRj8dCL+zeT+ErCh
ty2vDnnRK3O7tEOgkHDx4B3f7f7xRPUTp4mrr0HYezmuuBKT/B53u0oWF2O5hMjX
9eUEfQwjVWIBexVYp7/3gYmVP+ib/27fb194m8Eu5ug9nUnf8OAT1qpRkzL42t50
imLcbSsSeFIk80LVmBQ95QUUC912cymSBdI4V7w64Q5rFiChNZvcn4CCS82qeFLy
JF3Wb1dPuY+Pm3IOOlWPYQgxkIcqxjpR9XthkXw/B6DukmqjYWQQxrGNwhd0rwo+
UxJpkpCUmArNaFASENioA90Gkj/Sj7U9Smqr4UUKh5lybotxcDKXXTec3oZrFQ6l
0rSfLOVJ12mXioZaJwLaJUIW9G5BSWOgTCa+8YsDh9TgODRSjbWfkRuoR1OjTxLJ
3ptlgRA7fu2tv3zS8UTPQyiaQrtJ3ABF0and+ZbDRbre42Wr5q4k3enki1RplQm+
zldSEaE/gVloJHUSBx151NVJMFDtsLPS3fgoDnaX3LqdELiQ8Vpp00YCckt0xMxc
RXlpJ/hNAVW71faxNi9kIwrLnOYJyBRfYXsLJSQRI2wXWfp0Sx2iAucYigb75q/U
+8OWmq5vCFbdXRB3eo1PUuYOaXXa1GT2anTUdKqMk6XU+WyWRz1Y6gYn9KJ+W02h
Cbmz4NPP/8WKr9nta9SV2IXN2xYkCZagrFGYnGnM3nXYafeGQI/cWN+2YVF9u6s5
yVjXj3CGRJFYjFkO2FfV5ped+ObyGQHThlQCmVneXetJ5Pgqanyc/lw6fI2T4c/U
17DkjsmMgAWoLALVmZu8Rfll/Fig21Sa/CNiDdgAyHWqahXhMIN65GCa5d49PAeY
P3Rai7MzYG/4xaBJ1fSIvnfROoe5H5A+CZovUTJfWWKJmbI4c4WY+yliCY75VYdI
DfUaMBAHH6dG1CRjQXtj6y29wrrmYPmUY2re+4s2dZjSswRlwJZuovsv3tAKzP4y
4NWgH+/QV+SL6et5u0KvUDBCuL6wLYYj9Ig+og62kzXK+xkIu3KhMJvmqvpchBVm
kdRfqMWYOyXptaotJ4swo3TpXNiG8wJ3cXcfbRh0BTAhBZ8kCT+DhOOyv4NbvfMG
Kd/h6QyPcpewT2xPsZL1pS2emmI1a8CLJvII+LbTq4bzt5FiO5HH0cbRVsvFk+HA
7ArYj2grur7taCEQZzxUjVenAPJBqRB2JmrhllK3AESGVaAJw326uYbjjblv8dab
FzccBlEgqCrm5RixMq+V2sqtGyic0ubjbJ/Vbcjn+eKnxpiW/wc4YHV+7d2FFhUJ
x3syb+5bxIsYyYiFcE5v+zHe4cjVLpsh3xhBFt56TI/ST0fpuoxY1k9Img4MGdP1
RzYlKtYk1TXTrccBUW+Nvb65uAEFlRur62hKI6rA765T0QveYtUgvQEFeVqa4z50
cNw4RsAOSdvFHvC12LLXXiOzkGrR8G9CYXvNoapl8cEtWTFbwse0BGWTnCwjLSat
oQOSUSiF4n1+7Z/xrMKEjnGNG+jCbtL/nkH6GlglvSeq39XNhayo5xDgNAxwVm8K
hLmhgNLJ/YPGtEGGo2GyAdOXZTvp8jTikldw30Y2EboZKnIapLlYtP9NMVWJS6NM
SmpEP4o897GtlPM8d0woyiOZHSGehFpe66XZNfGkGQG0Mjg9VansM7zqaLD6VkF8
hYRCM2K9XOLUR+qOCvlBylJKZZ6ZKYBJVHsynaEl6hjiRaKKvAa0Vw11YjGRu6M1
2dtuzIdfm2nqQPrAckLAuYNRkHA0B6gETihFgeYrA9nDOH4UzvHgk2Srv4JJnf8i
fee28LGJjL6Z1hftTLmw/AOJDVaHGvlrRC97YTTmnxtGprD2aWDbxWvKnLGyrWF0
jN9yf/z4pF30/eMPzXrQwJQqUBI9i1mn/lJQuVHT0541gzlA2K3DKDRw9m3qQQsz
+I053bTpiC4UE9HI8uzNmovl9RG3wcB8iQ429eWRxm4Y0//8NcVRmyZWFnMX0kk5
5mMeQOKT9Cl38ZgT7ZPgHLsccDkiNE9+rNUVtVxdiatpp26TC9U/+wV0yG1NtAd8
B5CqKqupvoPkKBu0/0cXms8nkOUVK0U8Bo8BLql+UBEU6nXV4ogfziuZ1YSpc8nb
7Ad4lsgGCb5/AEeQBy4JYMm4A4bibC7cGa5bGkbeaVGZMPC9l08pQikrM7FnYm1e
xkg8/uX7VgMuMY4iyUKrIOdbacSy+ISSP7eXqgj3hmug4raWQ+8fSYYlCPI6nZGA
wnoo/6Z+N3UFXQP1wzF+l48KToRs2vAVm46Wcs5p2Bd9pN0F2CUs5vcZrhEAqZaN
U4W7ycwPJ8X2t4QV22Uq3Vr0Y0o6NBI3vGI/AxhFXRKLJ82HtQB0ftzoqROWWWcz
clbLeTrC10pbA6cwIjEFjEXdWOAgx8dXpP2PiwGsLhTbzfOuVO4FBleZNvqMxoSh
ZMFYQfyj9NS01ef0nBqjql5b82wlsQXDGlG1AtU/SDG+FWKeKGtyLfiLDjAVqow/
inEstsCeYcqEg5iaWaVam8ok5PoCUk3ZyuNSFTD8IoCw+yC3tQwtGOS3ZV951QUm
mYtJP5Is3MsN6f2wlp7ceCuOSAZJg/wqv4a4kZl4Z4pB0URJ8tbAYE1kVSl4qHDw
xdeEdzEFEH5jbLFqe/zj9XabRKXggIPpkeMQj+hq5W10MNTKdH2JhNl5C/yrmi7l
I22TP10zZfEt50W6ogwC3jYiBE7unYn6NMeSf4k/OTyHC2H6JSzWC83xYivtwN2M
HvXxwQxsw1nwaV46g4x/9ktdhBF4VawoY5VzO/gdgXeeIxQasWCCa80tGJs5Um4L
a0JN7lIGFMy8MylaU60nZxltYkhwqnlgxwAJZaEkX8Nb8y4SKPe6a14UaX4cakyS
+SwG+fjFjA+eBfdy8qDQSKA5FRqJvulEX1KIIhTeFTYagrxWR/XsFc89sjDXOvfz
a+otQNgUuMlLPiz1xyM5PX26yriVZgtwnwOMxq84w9fVSG/HCzDS5wlRRU+kCzTl
tyBB9dzR7osxnQSSYiY0oMoWiTk255y11jmh5s1nGOFM8tXKTRbaWovY2aec9qas
10lp/QaquV+s4PHe4ntbzD85uKIVpGDVNiHfVqFjBWnYDjlLGaHtuFgw9Sk47s+I
LwbsHuDt132ZNwzuWMwr7mX0dak/bCJ62oNJAZAdmqgR4adF6gfcKI7UbdJ+9lwJ
6qK6n8JQRIJGqeYAx3p1f1GHU5j2xxLNmaRUdESvMic2z3YmqW4dcVkEhOKYjKiM
v0QJHcS5Y/i8ITDFAJuRGHSNncYSooh79JhNO6ohf0RnsFiG53YENGx7vSLyMzGo
KHgGFDFfVnFmT1kYqW4ZDZJTnbgOIac20x9H8mxWc0eTEj53D+YrAqXFkQXH+UEe
lRwEs22ln3DYLHgsEnilC3sZ8HBglFga3bK4lvn2dB/uoSgGf/PchCTHe93CZfC3
aMbxpqKB1JFuNS1sYIWrhK67MIf5ZypzIcUUwj1ODy1mbbT+8BINvbC03u7Guk4H
Smr3YiumpzlQyTpNBnpzHPR3/7z/e0Vbbi0S40DzgvVe808QQGMGq/8PdBVCuLEr
vgoY7vpYxQoRFGRDOeCFj46H8g4OlzaNAgyBNfgZB5faFYq2C4ZN3S3L3btjq7/5
6EwN8UGxbW/jrQxUhSTvZPFoLtlz/WhwHGid+tFF7rmqn7pXRUaUJaasfJovUkBb
mo80JFHqgY7VQItN1q8zHK1CGnmWKIriKv7hhfMhZvTgOxSFi+K1mdRmqzMQja0H
TOpHX4eEGykq3DEiJ3/oeR6pGVcjEdlA2ovQA8mGH90gqIFO4Ed0KdLdjk7wLin6
DgrM6lHmOqVj0ByxbcvQIp+Gen9km2OI/5O5k0bSws5cP7YdYVNUp2tFg1lHZSfa
dTqD3455OLbyTyWK6iOqlHJRBph8ddJZYTXhPoFnkJKF8CmlOSVyezL0JdLmYd+W
BTrlkX9k63sTjNM2vRsfMdnATP0AjGWU0zSDm1K5qSEYvNmeoHoYe6OyrJI2Kr09
8IbTduQx5OG0D1JSywRjk47gAI4YRgKrDBXbBHlA7Wqefe3t+99LAdxpvi8XbrH5
NEtQCqwuWq3VNNb1nrmkmBYcQ43Bok7Az1E4nGBc6PVIGbSWSI5yPmsK7cPpRJoZ
HVY/H8u3iu7k9lXj0LoDss80n9THIqzGy9PvZ2mw1MAlO3A47BS96UHXNJ6oI0BS
kOu7OKPBtgQrl5tnMjqoZ6i0kEgra6/pc5rcayatQTRTMcoLPu+ly6bTeq0jcy3K
d8LaLzpQ/AiZT0nes+tbGSMJS9AhPpQMy4gtFpZGHyB2oB/M7f+GN0sGOUL4sjf5
AD9Qdd8TpAxw1cCgqFCRfdt9jVLhr6eqsWCwnEM1zxLAJjAGHXkSNpeniwuKL11P
kJ/Zo53Q7MibLfHfjiISlhy2t/unNp5ju2DHjdGZhiWJ8ZKDXfNr+Co5w26z090x
y/WUt/2Py7h3vR4sNBAvaum0KlSnU+zG4xVKA8mJ1plHDogXDWZX4bt5c6m82qk2
v2DIekeLYf6JqqTYHgdbBtHiUveFrX5Q43K03ieyPOPdfTJitaDAIo0RHOI2oKPd
+rK7gON259CJDCy+rsQDQ+HDREB6bK81X9+RLNRiPTtkmu/fMdN9FEWioWUQu3bw
iIE8y2AQdEaUUCmm5SJsF2/ETQhzuLvLHmJk+W4dFsMBA/dNZHS75hkubML+GMS8
sCaeMtNB+wtPgk7DEXYwHgfzuGJNxcqVWjO9GMnkpUkkwAUYvBv/Yj7TW2wlIFi2
gkGzbrlVuX+l4/hLNBnIz6ht/Fn3x5t32/8c7Xy90sda+cdH7kX5AJX3URR/wcCV
RU/M2irRxM799mmT+vcwXTevai46Ynue2iSpACAAKwb5R+5j2RFk1+3ejXw0FPyL
rfkTZzTfmV7VeOloY/NssJxQgHuGH5/qEU+EllGk1WfFsQXw/+HAlvZAeyuR/Y6e
Tgksg/6KyL7vuHaIW7Q2D+s66vpg6vMUeQa2ZcoyFlMEJP7c5cXbBAT0cqJ/zrt3
k06ALIpuFpIEcpgF0zrKi4I5Q7pIZknEdUEDddbO+awCyBzvtqRSm9SKuXrdBuFy
DwL6dfwzDE4eHxCn9Qun0pOXOxywCcTbj+Iv+TJ0mJfW7gNaODq76efIDGyuLLek
0PAts5FVgUHK07N16hsNXQFo6nbH+TnqA8czfcAMOuhUM7tVbHwQy0FlUpMhE7/u
095uhPxah82tniPlF/IlIMv7e2ER4LjiSyMmLjnoQpb6Y+kpYixJUdaBTnFApPsG
nwtL6vpLdQrGJZ4K7tR5SnS1yXMHqxA1ShJuflYNxI62NW8q4XOq/IDBmrursHKA
8w6fJgNKzdPznTrZca41SIyCMu7Xzu/TlAvgF62p3Ksdg4CvM1PzIfLYHFWDk8Jv
wwk+nK4TgVhy5BRqrr6vs+EMnbMKNsHE7rPmDbXyC2Azvx69J9kLYHewsgFhRfgd
v58XX0IfJP4uX8KkqlbtXq8p1J/XN+xkkmSPOcjECeFLkFj6R+Qp5MSSmmN0cDpI
6ydIQA8fRwkercub7dci3O5lKv/MxGbfm1GOhaqxUttloLsdpyscr8WmlxkcCC1S
p1hEwsUmQvVyYntLXbf1p2D0UE4gI8deZBLkiPXv1ni8NK5V1Lf25WjWkckjJ8HK
1WA9HZaDWgowET9ptiwDna4yN+SbAcUWpj40hB5cBqlDC55uRll9gzt2UhqhwOWW
Yox83naN1WLSuTZYD1H7WGJRZsPOqr7P88v8J3twQUabr28xo3hz/6lMlVkupJ5J
m/HWbZp6cRC84+BnSh86znhszWE+z23bCSzIVwsFuo5yBazvE0hk3Rhor9DWyN38
zGkRgDvGA8kcwm/spuNWXikHD/nOePgy5PsFhMEymVn0Rhtq8HkwM9M4CmvWtCsO
W5xvrNka1InvZ79XIFq3TJoW5+69qnfyWc60V4Xx/qDUTTbTJr8pIKnyzWT+1jLd
eGVXmbk/iPAUeQRSA0L4IPFVRjRU1PMLMJIK9GA5kioBzjHHQkbdHStIgYgqzwNd
8hvB5ICga1BrnF5unBLASvtfJ88vcaEV+oXHKN1M7zY=
`protect END_PROTECTED
