`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrSXgGkXBmErxUjld2kyXfiU7GaReJ8/kPtY9SgSNN/KGG7k90aJyDp3cWd4M9sm
rqShmCJp4WMrqm66pgQo7WQpN11l9qAb4uenLRb+/xkaqupmTs+6WQhLlwHp8Zlz
Ihg3jf9dgLHpNo06rOwcu0EEcaaJHau+odcWIMfhjUvkvczpeNgCKSEiIqjRf8cD
KsDzptSac189/jn3F4tCBf19+PTVK+NFXyHxz5VkfpREJbD99GuES95duGVMQT2G
sfAFNySqDyrFt8lS1+hShAe7B0HS473dAv9cQ8Sw3XW5IGYKq6NN+O3NVRaXzbNZ
eTmvvbFSUJp1aqcXsf3MW5PXBjRzRjSu9Pzja0FML0GXSh5SXYvK69i1QeVEJ3/g
AocbGJn+LUqbPjNA+Bm7LgSx2vWN17SAwiJvpv9Ti8sb6YuqccoPQXrh+BbalYZ0
DZFxXqz9/PCJ/KG02PSH+qWxYWX3tGWQYr4VrgHywuqJQMJxyHfh0z3DvKmxoomX
0NCDHfPl56DkB02mkvrCc/YhKpTkw31/2vKiSAQhvHaGXTRJbjvrlYs3fMhdiDlU
e6iyEBF+zFWOMMbS27zVVQrvh5STus5ri+7E4oTvoCT4sgP4kv3VpySRNCrlUXa1
tVUVT1J/mVW/HxBXjbN5PUSQ3gDuxUJu1Acup7mTrP9kWg05zhrtbt19sdTk43WD
avPKU6nTdX5iE22dx1YVFTfzGu+yo98GJEvA+sMXY0rZYXnaFlps2Q6mE7X6NJkn
a+drER2lt1ZkGk+hVWsqDizA6kf+T2RadFM0yGSq9xNekISnv1xvGaVw3mH7rJwo
IeyatAxeu3NnI0fLWwKE0HRqboAIJNFwtgKNptPaKBn1Do6n9aPIPDOTLNNjqeUi
TV7PuicHNWgiKKInvaI8IROFNUGZTTLKOfJeMKqIoI6vu6It287a1YwF2pnBnhFJ
E5vrhOXgTtAi2UyvVK5DWAlf1LE3occWal7vYPiXJ0RlecmMy9Rm27lvmbTSvGES
WIWIxHorpiya+7mcYnyzkdGuQliAi5QaEs32WNOkjrv8vchdXwyQcuXrXE5jTvk4
xxAoKLx389vtQuv9wdYN+sZ3gcce9ofrngqH8V+uOjj5ElpolFiAfdATaplFxBV/
SdLWz5y+kSaDpmRuRiEOrEYaiu/BNszq8ogyooFMSa0WhG4xpGH/Ny4iV5WNNcAu
gqkEYWwUO3tudM1Ce3HX54rABP+o7F0AL8po3QzPmFeJ5rumrR7/XyASnqa1W82y
C3HBgsg2PvSqQjCIafNI+6W/pQsPlh0FkHLLfdsORgXV6HbbmpJnafscFWoPoUdw
4qXpxOEthTMV8+9me2i2gteneyojn1pFQeFMY79GlOrfeWwGtueatCQxpWeCiVLa
yarOl+fkXlG4DX+kaXlOI+l1QmCb+k+R3qbm9ydxBdTYNPUQ/iBSzLH8znPKh+hQ
1hc2Bnz3v46/61NRJZP7/h8LP9ZT7Tz9PBDGiGlExVWNq2IdtuJE+9VUen+DzyEr
wdpbKtf53ETKXR6aDRySpri/c11uI3AN0TKUwWF1P5dXuYxUcQBqkW/7grFhsL/o
mSvvaNjsh4Iui4KC0kzl1lMXFHhy1IDtYEFyXk3+q1KWcq9kFU2+AuxJsFx8TTOP
g/kkeYLFteFgMRkhBzZIJICjyaEKajuEKJwG0AHHQFUFdrBN+godUF/qK7qSe5sZ
z0/yudwQIrSsvNU4oeiruBJ4TVS8PNtvn6grHOgbBQb6xJAcK1n4BzTB2+wD0fa1
QdpSiTfwzd1YULFso919au6G9iRjeyLDmtzSvANmALTiN9MkC1qQTYUoV0n0eXVv
JvNvMEgRUiCvo/MxocSXnwDqi8rUbHd/bqStsrLh9B+NNYpIGlbztXx9U8IPxNkh
7fZFx5W5xxH2XROg5Yos2LSKynzKVRRNO1Ky2GJEZ7RXA8Iyk17rDCBuUi5BdP20
S5PPKlXKSyVhBJ9Blte0TYet7nz84/Jjggl4A8pj6SQhSbOHQmZc/GRU8Jo5RSPq
nPDnc7cMwgdXmlc6wxelnySBVhv5o/JFqSxMtJMqfsH7MaODEdfiQHtE/gSWpUoI
cAdokXKFeSCtRsxF1HhiJ1BorOEudsfM1H5gkkVPcaVvsa/CisQ+p84OCktEjjpO
pIeL4UnB0suw6KYHPD6SvZKZ0ZtoiVEadQg+E3MT817opaitl940gOgfM7/hIcRD
V5zfdzZTCZ3aY7NoyFD3eQ==
`protect END_PROTECTED
