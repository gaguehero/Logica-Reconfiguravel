`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7I59l6dgEP1+aDUErV9ZrOvsFRz0Y+x+FvhkrBbsEfo5CpNvfc94UNfteMp04OYK
M2+YPmj9Uqsrn3VFrgW9DLQQCrxFgwvYpT61d65GXKtYJBrw6gYgJYHEjdn1a8Qy
Q+M1Y60nhOuf7MA3Mgw4LFzXzgdy8TGBSRW/e2IerAtaUuFEaRJtSoDVXAj5eryS
U7g3oDzmnHafayiEv76gMg3bzy/9CthpqCyO+gsR17McHOWXKqDrsFGCdxBuoNey
O0jCHn8hj4dTlDu4kJKUIGJslIK+RabF+VaR2G2IgWCIe5EvMz0f6+I/IpBbMXty
gGcQSAaWAj/u4SZqjh/3Ah+kjltosuIGEFBjvqyw7QTBUSulmcrBgvnDh0RV2puc
nFroSASP6H070wej4xZ6AduRyRKDdcaert4uwYN/tGXIWI7GyMFDDFuDuMAgtYuN
8V/qbE43Wug2nhWehhCUlaAcWBuPIxbzKjA2eoher1BunzReA78CtNnVN8BiU5YQ
qaKNCyC9YsIu6iCQ4i1RuXkZz9rv2AGW073YVkDZ0UNCAYtno/S78ja5yv6SRuE7
7F0HmKKQjytrV/meJZf1r2+Y4zYBZmdOqW3AgTRcUFZL444Ka/A5flZl+Sm5b6wC
x1qdTSw2/Bkb4Af3fvxrM93tarAxd/eHUc4MiO4fV1rBu96OTmYl8bvSVnqpVT3E
wYFevfIA/R/PajF8DXvzrY6r8HszWpBAZPNa/uRDAuFggcwyc73OonqszxSIpUFc
GEaGCZ5eteSAmE3BdOcnVbuz8FBcJjXeHQmQ2AT0gqJ+QBdA1q/q6HCMKsHMd1J+
BFBtXJLTGrHKQBLL8KBVu9WTLIK9mG0XdI/F05x2+zPb5eTftpt8elTbW3HS5ird
s18T+qQ3Qiv2chT1uWR38vHRoJ7nKsE2N9q96f9B5X+F+oBaiys+6i54XUnlnUwB
NhXF6gCBtin1YwkfWUgbNOtyB7HLnO9KNrezNxbeU4jgAWZRjosun7Qm607vn9/A
CnQxVOFXp49+5/4Hir00KuRUbHvJ4bPH8i85MK1edCpJWrmD8nYu0LPrmQBw1AM/
2ZIdfzWfqV1ydGygMfA6bWSq+I83SI0Kfoo/fZZJfseVFaypgzBf9onKiWulUJnE
52Xshe+mddM3dk2Hnmq/YqDjPzVQjrhf+13jrVzs3jBH2/RgMWPIvXepF6ZyaFcq
Nzly3cMvHK/W+WNFn9ncFuvlXJFpIs1hxcFcbQGoDwHtupn1DHI98VrObTcTz7Gr
kyQH7kZzlhs/4h/YQLRS7uZfKiMnFR8omd9V8D22olmmym65JvcU2HKdUtQ5giK6
d1/tM9k8TDSXYjXJ7+4lTHRbMT9q40SR6Ktc9AbwRFwB7nfWY5Hm9SSaGujct9S9
2MZXQ06VSdiS4HmFz1pSDFL7YC//xQfwp2pY0Gexvk2pWViMNSqJlZxL7zmQ34qx
EWg6OVCMbqfy1Xor50v1CKUguR6nQ6/cLRZlwIGEGKfh/B06KFcQjTNmUtA+Gd07
50KNn1tcIqda+J1ioHMcU0xDDx0A6LmPJwWnw08nwrT5TeWJP0XtzprrgrGVz29B
oT4gc4GkhEweGbWEvjD9KVzRFXlN3Wf5sa4zuZ0SKzF3oJM/yJuLtlAXnXeORFGH
+VSxnFy4V1MTg94w5dIx+GaPqoPBW/ZV6lIFTyJ82wLOAZVyD7WbiqKZOv3g6tYe
4ff3Fyvls5tdMo0pUARxpic6vtWFrSsiTPTrXgTfQ/C73A5tVtyn2QuS91PNHXVp
Ag9zK0QpUgDyRIqYbXHlFSDiS6U2jYW+qznnuImshpXYD9nPzvLDqcUyNFDmmgon
BJVpr8Q2qxM0Fy5Css5NqjecerCkdDuGcFO0B1sMu0r3bysiwYl2hyqjzWjoy8De
0KI8Nh9z/TfjNF/GiaeHUbKwwIrriyc3TIxnNY6kBGOBIo3rCYfvWe3fMW3wVbKA
UX23QO4VbcVBZMCPdn/mSNMh+yea318ZYl4LyH5oOHD8Ak9H8y78O/yjTVwqSI8K
`protect END_PROTECTED
