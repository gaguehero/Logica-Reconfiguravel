`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBdiO6D4yDvbk3Y+d+Bm31ihqkwRFHtLYB/ypypHX7Za0CZfsXC1cHaGSF8Lm8cQ
JIXQfHuKBe5imZxk94Ru8NZ4TFTpK4poFhz0avMD2/uMMAjXyMlAn/r3su4GLHgZ
noR0BEdySbC9UBf8KO1XgxKmuYWAZH38Bk+inF1CHWX5Yk6jADjj9t5cTxJXyiD3
zdoWOXhLBySaHCHIv/n+31kKlYKSJgkz8t2hLC3tyvz7u2ZXcQC1gIeSmHQ7c7QG
c/z5J12A/AKQSTIrtAjoDQtQbeVKpMspTGsABR8KaFoG3vlA5QJjYaTKKYAvLUIl
V96RMKSq06OuZbwbrghinRp1aalj3VKPHrTjG4V4TsoFs70cHW+R3pdG3I4tZhH6
v9z0kQPXxFYrnFh1ax8MjZ9mu+fCagVJbWKhRCr7CHQFZKu4fOKAGiZkP4nKSb4D
Bib7BCaAKNabXDq2nwigiHKWG3L1eQVbKd1I3Fuo+yKpnSkvVHntOYsVEWVNB0Wa
g/D1/G3APJNH91iRxSuWnt59+fhgg0rOQb+Gx4lWaPb+bNw6et1ArHBWn39DIe6G
xOCIk3vlYyEcGLUOVawhaEhgOHXmf9n9GAq1IUiGeqrFDhYxbQ4Y1bRVdkp+XT3m
82j/jfVL+TWLyNzWxMGzW7Aimj/HwFXow7jCfCDmXFNa27wgaaOmkClbQxf79AOQ
+/VA3tP6xPKsE3VC04VM32ba/+mkgGSGID0rFV0H5jqy9YXRYpyJsj59iDuXnMXS
KSw1lwbSaHnAfy3A4JP3rN4nRu/RsHNrAX+9v2M/jRms7E2eVHyrCkCu6VlD+ML0
SE6zFuCITbmMblUJIBjqkRDbbGclo+devRIGIbvRkeOA1qmnkX1fOIV8QBMk4sUJ
Y1SM0D8IhUaicIzFMr6RiYcVqH6KbXjJ9Abl/H91OmClr50Gxw+boKZ9Xc9Ex3yy
GW4BG020TCjCasGFui1fS/QKahZyHskH6i1SzpnAcd3b5o1aKRN6GnE7aY57vVuR
ivOIBjs2h4gsMl8hPuzhMpzvH/bhz4ZkxkWHWymS7/gyEFkqiar/6UncpsMzi3px
GuSxwXaXH4qG/C9c2sBGsbxTku/2dBG1tsX6sgG8Ar0E/QqhZ6ruuCcnvMUwyPDk
220OxoXEcyUoXNs6OXsqTJ6vuOxPPNLa6vfh6ozO1pw2RvYXeT5HK6YpqeGRHqS4
yUurZq0u+wUIX++RxoKY82vYQnbfACIiU3enj6X9I3+gGHVJtPb8zk12gCQc/x3u
NL1tzoRiOPGqt7m0Uwn6GXaghU4Acj7nQAUjQUbDEWLIJi7zwhlRWZ9cJEAF+iBG
RNHCIuRqLwX5rH1x/5iMYavCc+LsdAv2VlZDbycmCfrOxJEKjlsLZXnRJ/wA//ju
yg0VlKfxug08TP3DJbBwMUos/8M1yfijPRrL5TADh0XttX6kYBHOinOBIwlWF3ul
ugbPP0WHEXVz5kBCFTOUohP46NBXxQA3kFcmUp5uD8LmcE1OqMxZO7O+EA/w4GED
5nzyk3PDYRay6Z5siA3afuELWNnP0JOQPj3RJs2uR/yKl3PKgtH0h/9CT6gND98u
GhuAnM2Ev7wq96lUqLcgGJr6r1+JLkG+nMNpas+F24KR3j3ycBOCDL3HN/iT1bBO
l9MewFYUQoAFA8WvPntUnieO2+YSHrHz1Hm3x126l17Hiysr24R/d0YJ7Cn7T31e
GGU1qo4RqU65vLYsuZLsRjj4JuwVxwj+eX1lBsYFUyRmrIirYFOQw7tKh/V97Jm+
mOMx3ro7SHl9ymxmzvW9OCk0w38hdACwAkvSQEOK8Q0oovBSavMpxtYzfmq9xNFg
UlUxzow0y4QHMS7iBDSOPH4LprtGMk4GIRoJBa4Zo2xUyaA0O+8P6phlHXhSywOn
FhtI8AXBVl7yW6EwyMPWavX33DESGOShWZL122F+8z/JGTmoewF5J5at94gmz3Q/
OnD2Gbb+M8Jdqs7C5KzbGbreco/Ajrr2Ztr6MPQDiWkMsDECFKFMDLtp8BBz8xNo
SWXYZar466s60mVpbn3IRA==
`protect END_PROTECTED
