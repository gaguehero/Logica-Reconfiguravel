`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BQVQcmISrss/dWC+Xjg15isFV6dE8sn/gYXmmL3sOOBcaZ2jVvbVMvkI4GvpHxW8
JW91mwxqq03ypNkf6PfeEcGVKbULeXf8gSQuXoEqBWPKUeyAhHJCix7nyrqBNPDj
mOyQv4RbD0d3KgQVe2w6jDHJPYGgpksJ0Vt1y0xDHneANXBy783KC24sknlpXKh1
p1vFPEyt1Kxi5ri7/ytx6TzqBWu2RQ/B/MStGNweVczRCaDm3FjM6rYYKJ3ntuXX
7fIE51RK7JRhD3YcxaOpOKsjMZpT3argkNPZn2TOfQFHkWQ4CE0/5CjBnz5Fm6Bm
cVPAbP+zEiXwSP+ujygKdctVgk3YHC2qvwtAfKow3OvbPpfp/t2MR8bzUghy8bx2
6hefPZwurYM+97LmxFVg06sYLMgqllUSigGLIWjjVAZIzvYso/SJhRNjVJrlk9MS
/XbSTY4UAjZbkiZ7HtFrBMuO6y8u73YRI4whqz7GPPR71cUWy/M2c88QIar1auHi
b3K7asxCDo33tbj7EbYQQeIOZBo4RSOG8qOWdQEKPnzBlYT1cDU2siiyrLgBinqe
SmmrtYu6FAYPA4EdZ1dsSv/ImKEtnFvDNZQdkqw23a7bLtX+IuN9gLedp8rKy1jz
ZUjCMKTbfahWwnvwXanaC4EmlsmHz/ABeJhilzPEFG1iFlp5IFJUkaBVFHwVUXZm
Lm8CEJzrpAXW/h8uQWJU6gYEF0TZT2lBsh3g1FS7rRQhp/L0w4cQdr3Pe2UUqeuk
kgdtX/N9gc/HILFH3Dk2wW/5k+BtG5jRgFBSMXAdnj5dgOzs1VcmlCKR4g917Cwb
bUBk+jlBfZL6jn3J1R++FTWMAay3/H3OPRu3AiFxK6nCY4Oz6UfkFFEO0gg2/fUJ
vLznYrAJ+5mTmynszHYSMvnJUPlx8xi6a4n7MwvTAx2+8ci7QqY6y1Np5ea3q26L
kzw/xlHlJBUxejRA0SlkZ5k0/elr2BD/lYtIfEvzEsdlmd7ySMeqlRh6s7FwR0yK
d2r1X/4bAl/ZrzugR1uVAXUri20yrCvlFG9axB2qTT9xXfdV7Y1MCZg3PXTKDRFH
AnMYc8XFdu+eXLWf1PYzpfTphfU+tbJ7bjTc+JxN0j8oWHmsF5CkwsZQbiqh9JQf
Fe2SiO5VXaDzZdrP1VJYyGpzLL/xJzsT12QxQ8cxLYxesN7Vvj4bP6/v2l/0ZniI
jRJ8PACwOuzhhnnIDX4sFOlONaLOf8eo+UXn6avA8NINen4dNp/gTXbHF9QpEMZd
8e+jUwPlEj8qhjTdXqr1gyA0ijkHMLv47Pfnq4ZO3jIqSB10M3UDOp2vCKT1aaav
ZXDtm1PTRLaVICehS6Wvud4uExVo5SAtXbZtxAVBPmrFx5w6rpB7eqXGxKroQiF/
2PosdOwTaMA5mQkF8as5VmorDUvYzQrI9zALcNPBpAboElf9ddU57NQswA6YAhZJ
z2sV78CmI4MOhIg7KmVFJbeSCSejG1e2FJsmt6F5io+7lO/xTYPPLXotA+JuYB0Z
3MJVVesBo/B/qwAncALZyswiQ8oTtDeVHmGW0piOBlHy3yDokBzEvxNC3agkxanh
7NBGQHU18gRUCOoOBaewvxxK5doQgu9wUz4fjCIvYjEPadPAhUSoenWu7dMPfYV0
P+4xWIOTzmH0v60+fv9s46vvDMn26H25tqUu62mRnAMSECaxYdv+DhGlhbdNPtI7
oG7e1/WnzlV4iVBhfwMsW44xl60xMAefh0ei9vijfvEEXjWNY62Lk7IcgDJzekh7
fw+VVNr+dmFhUqLhu2/gVVGAduPqcImpZ3TJ5PdukQdajy6YcAJTwKDn4eJ5H6N/
CFNbwKv+9Gza7UjpS3ORARC11VDiFJzn6hwDUctxL36hvd7KqPUzExHe9Q2OZ4VK
z6rzrzk+C1B9B+FWD/GhlG8KPf/i5DTlEngiFgbIbfGU4NM/Tha/5E/bLQQwNYk5
Ghs3nyYkZK43Gxq/9RkorhZzjPMcSq89pmjnG11+sPtjsPTUj2GZnjSsdSQ0ucyz
n2F7NmirT6I38yw38DIqKJvQZ55wDJzEnZqjMIBqqjNJCYKO0HeB9X9wq2OO6Qpq
XNNdBb2uyErSHogqWR1ovbq1NZtXQzTWF1bzpbAKmejRcx/R5KOYDipBXUpe46tO
xK71nhy8mPrUw3BC4JpdHNhIGdGqoVPUb17XHoN8Ort9/3kP2RIxDSlamYZ9ZiDu
BmLoxBekKZIZQZCIxHjoJvFOiZBateWYKHiv7RBgO5ih2qnWCd+FrQe9eWfQPvlg
/xm3ybNQMG/v4CKJhQXgiQdahqfT9mHiamAjYiYslGVw6jIOEs7Ss68pT9weX8W0
lpRijFouxJuD8o6vkl13O/Ckk72ECMbC6kXTgcwBOQPK2JXCL6zT50m8nQ657pTT
/odC2FeccBQJvyf2Wd/4/e/zOpLyn68pnsWPCxV2G7Lr3JHb87J61UVCDN1/FdT5
/bn4hh9t/97+jNIbABjx5WITvwKF0rQ913ARyGiuIawpAF16Jeu/eExBNTI9LHUV
6rT9Rv0N3aK+0fZQQaakKMzERfW8H455wY7D0OXj9c61pTBPAGAk4JIKihzzrbUZ
gZDpxvQYqTBWOKiEqPSdz/trKiFeqaoNnIJTfb3uaJiyoOJS05hwsnxSn95JJau7
3WghOyMFRd5vZiBJwZOV6JmB9Gsl8x8z9MrSfwhwTwzrfIvMpgt/z5ydfWGXMKzt
AO0/raTvyXqH3F9fxHgKidgbslyws+avw8U7B6YLhj/0Epx1Vl2nlfkw/tfxQXTF
t5U9bnss9OJADjr/lCTCXboJjTtkYxGXeGOCbvyMyfvO31/Z6RCFdEFcye6NKE8f
1ui0K2j0qycd77fybwGi9GxkAsx0U7mDBB5mtWrdCbyhcVxvdnjR9vWV4eMSAaAL
Tb1aZimuOMfvC5QCaDSXFM1T+ny7lB7Jf1/haCCAENv5mRAyb0RNhVEa54CQfSvz
N8WwO5rYj6462soSVxKV9jZdCgoJ24Qms7s+ZIlGTxLyeyY180/Ev6DAmrLPOsZB
lOTIF5GIwAWrNwYilpDlmdeODCjXLkqhyvdFTN2CXKOL0VqNpo/JtU0alQgIBdle
M+QK+ISEi341Jzxp64oy8nmCPdOkhyoJ6H0BMjDMz7eFB+CMyRI1AOzHYFJdjpIw
kW97YQ8ZLSjSkJwzVoIreWWmDt72Ejn0BWQVtAHZPlPSE8ppVeV+Ul6q1ronh1DC
VrtX6dxUl1Cly18EH5L5ZgIHIv05nPa16O3ExWSqwcQt6dsZwoMJSBwyEdvuk3l4
f40Mr02Bsrdda8xPnlcNY8jAm0DVkbUXH/K3sOD9eiDWqQ/2gInyOlPKTEJ4Ioa3
4UGiWU7N3Dg0G89/beQiPNP4IhJ8qvVx9L98HLy/fKjYddUm7/IuwKk5A3r++ovx
ubychlQzer8NDPxUSxBYEpi0R0/2pRU/nNOhPu7XhvDka5t7v4PDYS7wGG2kZoem
3Iet5UqZWXJrGzUOMEVYeBfaTzUVC4USmA8INWnUVnzYTwyuAWWoWLJ1/FDCVjkc
T/J1YJ+zpQVDNvPFqCjoHCj2OQJBENoszsIZfADCrrSahlCpDWA+FhQ2KeTt63OL
8G/BoYe16NmxNDHFqJMiGi747Ok00pqMItaFyDgYQFy4Lfqe/0TGl6dxYIqOOzjM
UhM7gVt8Wudsh0ljvBZakVor9NA8WrtScr+ipBENvHFHNa21kRkmTUH4MYtYpz0D
fAJpXljYnlxeUkpzma8QsPk5Ds26H5dtC1MjCbXDanio75UaibbfjrqeV/xQo5ch
gd6FygI6HLg7ps+V/mmBh9ZfaQZxrV0f5WEmqnD3zZCrnxTALEQjCbl3Hmc4u+oJ
Hthh/aZwmXrFChHfzwD3iBEJAlpnMz/+CIDLKi/qA+qt7ZH8qmHAP9ny29I4RnWk
aIKi6eCfZsgg/uducFWu6mziEPEKwQRRl3/AR4YfvFSBdk+s9dZOqiS9PrAqkBaV
anrJ0i7sZ5rwzKGlsXHajNjBYVQIrmJn38mPbyAZutfd9DUluMuCHs6APTIQ9QtU
4uJhkcTAEtpa9HnjpxOIc6EKot1AY4LVraR0JpTtsmr2TNWYUdngldoWR6BCtgHf
s/BqjrmjHUWwh6ZpOp9B6Du5T7SGcBa/jOE/C2TbM/7y1DfHTE+E9m9puNnKYxR5
GN0p/nO78BuD7fNNcbB4fEFL69kjCf0VWb5F8QgX8DcWEDb9mRBEJcyN1g3GdLuh
JzdMDU+5oT2sYnw11Z8jUXvr0rX77H6okz8O9JMIUOoHRjhNRs+au+YF1SAqBPRB
t2vKgIcpAIzpT93QByqMons/rKJGDGdUz94sXOUs5Ar8Ofkv1Jjod6QoZcLBIcQS
ItfOO1ttoXIcJ2WjBL+7oY+/cTOZIClDY2+ANIMudb02dxd8nPgvmw07MoHDaIea
1IQot/IJy+uSBY6ubXJ39RUnlFq7vjIgJAkvo/icu32Ou9Wq4m9Cib1J+t3xadUx
pbvaQNRYZaIJL5/fiJveblA9uGHgB+/4x0NXS0ZEUMMGuYdBeQlGqqXsJyBRKxe+
i/et9vC6oRS4VgiWS4oNYMI/5Zyfq8LxftWqRzuGW/pVvT/AhRa7gBjT5iugWofk
qvtmsalZrBCPWWBGUa4KhYaKdRCcVpBlSyqIsnISjXgAahfgg7gLCZFamiZBHdHC
KvApnNSHYscKp0uk4PAyEnFjMLWa5jvToXiKhMdMD+eAKdEO/LFflOVzQRqwA1Sx
Bas1SF8DfSiOjIFpPKU7BhvFO72/NAc6K7flHNinkq5t/RW2n6sud4FOFWuH+E4o
pcPd1DsWUKePYb88XDVyNg6BSqF9alXVGsozvq4F9uvLsMQtWtB0zZxxqChGwRVp
sTiSdDbR2RhmTP9Mo93zsqrs8ZsYxNonEqpulIu8gPdF3bNCCt2b7Tcyz9ArPU/Z
gbX8vPbg0ElOJkornp0aTlvjyCy+8oBjRjYwdy8T1DVRI6oUeq1GDgkfcepPVz4c
ehbpxg9tvlAprDvEV31CVLZt2/Frl8GeGvvBfi2tjVrs3H+dgVI66Z9PfBpe0zyo
fqV+capNNKS/RzZIRjfxK4WlCNj+HCzAihye0us6B0g/11OiI9ot9wPBq9Z4WPuz
XAN07e2HooI1Z+3JoQh/PrFZ9dY2gRe+39sV4oWrHHoSPqFavkKa1aFKoI/+xy1l
zUj5z53bY/UsMJ94U498pnjnoVbHPKWcYRpuTJ8yR7dv0A57IYZUIpwly3Xu6zVW
kVfCUu9IDma9E53MNY0eJz2jPspdasa9EwD+mobZMdwiwoZlJyH0sdms3XxLFLP6
oHXg6a0ZrS+SU800jpubNh2nOuCO9EshQLahWUI2vjemWGxlDXytbDLiVl+hewuA
QeksExpNoZo6ASZEIdbwI+bVM7jvvorwSEqATrVyFDXjl7FUs8r5xtPhWQdmM0Gi
AKYbv4GvdqwfUfyOBWmmyqTVWo6L4TuZEUfj8dOXAArBCTYpjOXaufRe6exXofOX
StHnXjgmY8AoYPTc5HNe3m4QrVAi3Wj3F0giZPAPAUz0zAF2XbYawmq9JAe//kkm
A3FaZCx8DraexAb5uDlpBCJ5ZJ/S88imS2tACjzglSxWk2efY6IPxIAbE8iUveWb
nu/y2/VT6QM9r+TgpBIf8Rc89oNchMftu6kvgrh0dqyXct6O4ngM6ZVZL17W0kHu
0hP9sToOk56nij03GY0FsXuGQaAz/wGBsnDkdAe0/fJsZqvPotBTsc6axnLUFrKK
pr2oMRz6NzyNvpXXELXXPTM8RQmH0f+uMbbEg/w88pUAWor0hNCnARiZUYO900Qf
rveia7+/RHCfy9djICZp30PFL6mp7PBtjSLN0v8LMC6WUQYECK5GI9huMdBFVs9V
q6g/MnI4tER1p24mkYUvsGcYOxvxK6XcnOZ/3K04lDmYJrtqCHXHyOMoaq3rAymp
OIlrJv9iDtgD2vcNx4/ZUQjqI4Ol0JtOz/PNxw9740K27xJmj43cBYSyYOy6xcI0
xB8KFw4kTZEkUWgxbTy5PORnqOBN7ikgU3FshfkO7BXNcKN6KPa34lFKUChTJADt
QFpwPOHiV2zPvW7PS3Vm3sFb11Z+eni8Box9N9THTlZm1bN+QqqtcZdDnSAeGcHZ
7cNAbxWWmqLtskksukrnzwG/6rVTEnJxouiMMzRzxkGoyd+6mPfG4nG+4Ba/wgFy
ll3gSpfU2AKIsEu/hcg0CK59/IFruzVz11MJJO07Rt7AEc+1Mtuh/ZlgFcOvsxu3
8mLPSzQl85PtTaUqDgcU6Ay3+lowGofkL3HyUs5O2tNLZzTnqPmWLZ5x/uFzoGTI
BFyTnV1SePbBnNb9v1AM9Qv/aVwVTlVSSVeVkMh0ZTRrfFnt5jhezTBbm3Xokoy6
dhhzC3hVA0yMcPw1MUtwjUQr4KCSENZMKFbHenbohJB/uanYWg2uOvsosijdur2M
nwyHdqp/pc9qs1Gefkbfds+mhVz4EUbq/yimQcjkOlnPHraCpfGD5P78dNlsTjAV
/8KVJt20+upAk+S5XXP04V0hksE+NotvCw+HyQ0/HPwC2zbtPJ26PNMz4tyvE+W6
Qw5Wvh4uz24YMaFcdwVZdol/e3SqQzPN0uvk3C54cMzJH442TeuVdQRaN6Ugat++
9pi1Hp2TVqNM+hvqXfh+0IPqkazSxX0lm4u6V/yo7zjeSoiAbWiXHmkrMCskkSjx
TeoXlBQaJoyoqaxS+dPeJUhspBbhaDHoqrg53iTxTRZVx+9OtJjp2Rs6CWh5rrvu
t+zRm1z5n9v8a0U+o5w5CC1T5v28NHALUV/dU+wLdVpdO3M2qWCYoX8wPulGcjPH
U3WVLoIPpDV8s6Eg0GnePZHLr6hva+q6FUMD5EbdAkrR/mp1y5Q33RZYhMZvRHzv
YCHdO8zqCg0HkKmvNefY6plVZs6LBBwmRLnazJQSnCIeQd96Cw+vfSYl1YRWnCST
CjFoH+p3so6GqG3Ykzc0u+2vCNxghkeN6TymM+l1U/ZxuZH+J3mghXpRksNWu4n0
enpI00NS46ST0KJ3DXg7ZrjX2ZVaZiBkCb+XsRS28gtPRFy+43ed5YDoJBx6Ip/l
NMYG/upyIZ50MrESK3NH8TtE1wkSXdzCMAiKZ3XyDlA59as2I/RNR+DcRU7+o/to
E6tICvYP65jLfyJWx/dCK2axKj7jWUwyEA3FmlZLDbu8ouHqq7EYfKNFGwwExkiz
MZKnyTyZFme5CWHNSfdrDVsWJMNJU5X3WKj+iLhAyVqTnklHzQ61j8XQfVLfD9S4
xdX8dc3DqIlM1Ryqg1YWuejPoShBa0wBy0Al7Kcck0zInWnr9tRnlX/Zg7NmhX+T
c+tsX4pZgqcW1BOSQGbgE8EGzPNPZ/8mV8PXUB7vhWTeEcjl702lcbLhx+WjmA/y
InQbiBBxf0sZeeWgW508j6izcqJA8AkuyNY29b+MoxjiOLiZYhyAGFwnGrnSXtu+
7ZYLBX8ZjdVtOKonDO0Bj0KE/wGFMx6uvNt++GHpQRl/0Ssm5fcSTZHYEzcyRPi8
BHF0TbW31yiDm5liH8s68ttfDgmvHw7nGci08fUaJudCiTs8cFZtrYwDAl2F7i88
`protect END_PROTECTED
