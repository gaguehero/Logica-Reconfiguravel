`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0w6KdEoQTydwOXd4skAy3SutsHmigKaYSUGGRQ83qLzrzbL/eDclj6s5Roa126gK
VPR1bkiPWOQFCmOveI7sXGq8sHbABcyz/AD2svBcM87vgvTZrRzvDyDGSLQTOHYe
qzUNh7NVf5quZ+0LrYRCeVQSSjb6HLjkvGhnqf3WYQGO5qi6Hu/jm9b8XVzO97uu
i1jlZBNg2bpaZdP1q5XZDKD4GkNJqB1pOwTl/p+eSJ3KSQ4s1S8ciaCF3g9zGgzm
wgn/PXlGl7cAqgaHb6bIEO/cZOEJuU1ejhNMbGyJGQZjUFzR6e6Kl3X2yAUTuHPf
rkNrXywjXbWYn0tAe1bJbtfz96z0B8v+0DPzTs7zrQqQ8UrsMI/RC1wY01PCbemg
GgJw5LZbxSrAZ80NjmTddyKFBKhvXZw59r+iL55H/KLScY3YG7Oo8tYQRFLDOTVr
8IVp+9H/CtbLlKx0Ab5P6UxddNX0OmrcmevmCbLB2x8si1JlrY5mTnaUhv+2V5BO
mrHLIhArBEvTSRdT9Yx3id8y9C82i9qbdLTcHM0/wly55bi7G9TU1SP/EI0FW37/
HUd0H5W5Dm4sTps1IwK0Zw7PbrNOhpLZYnOK+vSLHaR1H0ogeRokhsVZFIhtK+NT
0lebK1IWk4DhrKIAGFWeFhsqkgeSnMH0EurkQLwSFjJtv4sySF2BntiQ2jXx61P0
f9WfFE3znXDErDwiJpJCv4zgJIhdaQDJqtCnzHchEN3Q227I+O4K8u1ycdgmyzy8
ry3gFuxFcf6tty6mUsbt2/zwhm4bYQCnltnisEwpQRbCQHbAQALD5bnSfesIutRh
hJ22Q7Qe1jAJ+IGRZlV0XQmf8n20k/OA4l26vGlXRmag8iSV5xxDEPRGq3/ck0mV
O1djQXNIux+pmDWRhrtdYrWsSyWc17eA/eCfjhweRjttSP6Gt2/CpDm4xDU69vJK
oRJnuWCrtpHCvpimZCeFPDtDV7gCGFLhDAaYFstqnFZs1L1c9n8WVkbsfvfv3SM6
qH6JSEjeo0b8q6tHwXCOdy5RMIArJKdJGXt64ZVRz26xDSGWl1GWLBLdBOczqWiM
N/Phe5iYfgs06ozChHpUJGWWkAIsE0nyCpgsYEemE3X75OVN2o8vHqBwNM7Vpn1S
6DqO70uwlThGZkHFeSFvpLwxhue7YzcWJsuIJAcL//XMCnXDcvh1F5+i3sOV4C6u
zfqmx/gLAFWRR0+3RVg1REYiSlCBr+H5HiCjOyBOwYanGpYIqMnwGOYMqhWINUOe
vBXPRu71wou28h/n0vNvqSkTQPtK9FExz7YXx/b3Sp5mF8HWR+fzK39toc6dhURA
fNCt9kcZuqL/M3YI8fSBM/VIzU+3ZDW1jSil7rhjvixcWZ0UdjwD0Zx9CbpkuZtw
aNgXsL9QT6VQP0stznIltz0MS/ht/svMeG7XJIdtGKvKyZ1hfZvKrRqYPYNpLnOw
7VBtmbSTMimt6KpbfFxNYUNhN0skCikNnVJNExwgrEAVf013CMPHaaNYWDA+yq73
OmTceZAZRTwCvLtj60fHGppRwU1zEfkAeLUm/jwhItATmvfnYZkE+t7qWH9HUZB9
SIXa89QtrfOeefdeuIpNXGyNuVlW3T3KhMJ8vAQ2nO2fHyFAoER6gQcARXslBYR6
DADL5w+QzKHbvrIcMm+xaETBVpwyymQfj2MmbiOjUWF2F6lDQv//TqfziQ2kDs4/
8Si41Vl+J3QNhSUI5tiEnlnJ2hFvko4nQX2AsXsv89GeGa9ZxD3jFnd71i6mVCQn
G1QEpDMxmnsDuRRbiNbmpLlxe4UILEumE+aj3m1sRi7ehJ0R9yBpguf2j1uJw4EV
wUdHvVrblhGhO+iaHP65vKcz8pmU24FUb4WGUu+Aq+GXnu4miJtU8cfgwxrFLrdz
+oHp5rHbLnaI9Sm73GUc4a4Lp8Bktsv3zjIf7iyLQ+OcBZNoiZjJ1jbAzBYXs+VO
zamucEw6zDY11fHGAecdm7pAOY+JF2QoKWJSr1msh6/g2y+dpEjN+AqUDBB6TIuy
90EE7zkub+wuB9HKj8dinyriMLc5dh93ZUZ6Un5ADZ8YwJPqFLiNL0rpadqFIxvn
l+IuJnwr8oPN6C2eVC23aVmxgdV5RGZ/ChKUZmPOIq1MOw8Wn6GUTSOljwNJfaJB
0Ne6AnXHigb/UM6vFgomJJa1wXTfUweXtDMgul/iSoCJV9bOTi37V1dWLfLCSdTf
8bbgaWfA/lFtTlJ6kgRi+yPkhQc9PKGc/pUwMFQDUga87YwF1KJuCNqLhOR6x3gT
n3sB9lK4HHEMGvigaYsOudX7ayckSPS2ujjRpQDls/9z8cLEelKkpWrLdHaxapbE
qr6Uak/0Bb55buMsZWjdH1fzv9kZ0BseN28gPLzNUg+HvF/uCCJoQ5AzBxBqwfiS
K5InQVUICDizERJknUcKpud/fxYxZOv6+V8WjD1FzYsB09e9Uu7+43fU+nM9FNFy
q12XjBVxuaVASwUMysZwz0hwRGENBnpenrK7pCPRhSCxreW4UmifylO+ghGoMwzK
cb01SVLdXlt9p5omCYZhqwCgMbXYncCol/zQJN73KRuDkPiGUBWbELP47Tts/5FV
h5QJSXuoz1xWtEUB+ppl+GP/jPUECC9QjjockBtn2vREFpgQtAND90kWUdV5njtk
DHnXGJir1e1ekP9lQN1Rd8h8E8bo2k0hTvIURVKhdN8sjyeQjALUoEr7TRuPUyg9
wqZt/SXAGoEo0vHIpvFUtsDyUV9Hv0/AupQIikXEXfHSXldPz9Q4qH7+ZnFiCGxo
5yQH+/Ng4pKez3BARFvKdVC/+lM/XwGM94VFkJ5go7KPjIeapx5Hawz4VZcNZY/5
YFSQvdTK0aOUBKPk4AyHAqoQ+/fcPLK+kLTxaBS9ymeLHXXprgSRksqC3qpv813r
fuMH4EMguGqLFWv3kO/K5WyHGOWdweHWQBMD7rLwzkBy0Cww7jS9V72cy9O0awim
841M6UmBFbfdFkxRYp5q791O2yhPJUexjBCNGMgRs6YSNL0trKh4vsnla8NSOta5
RazIUf8bqsg0EG+SdW21GMxVGXJJ837ii+TLbJ9sWoPGEbKFqkpUX5iZ1LMKHUFi
jCZpSunWhbMZBe8LI13Nt3Uyj5t8+uLA8h5Uv68NfTUdKS+dupZ/y6tJoXWRZASe
8DWa+ySysedgSOLVShYjAjB77F/iysKgkfRX9c4K9UCzdFNPGEiakV3aN58MWKx4
0PDcH86oAVKpXucQhBWU9Z/CloO9WXpwAuJ0yRdmWyERyNdoAENZcNVdJQdXie5j
7tc0+pZS4NMTgE9+GjjV8c0FiHnkEmpFoW+QBadMibxAPMwIcvtR5bHf+pte7GAw
8rDeEkRL/ReTFzoAGBqJ0DiVcj4coYlAxLmd+JM5mA/1e8Y7TjGR3Opem0t+T1nN
9aN4iX3+RUf6QrptDMPELKmkJM2JRDM/eTCJlwxSZ8qT79uVazM55CXHJW1Vr7eu
SrTkiD8w8MD157mWIihBluxgXg7d4Cvhwp80n/KBsgxzrOGWWp8tgpUdmF+h49QF
WN7yb6kN4TaGES80Cr1bxfJlSVFtXpQpbWHnBQyxSwa/Z9AWpZ2t2GynSjIybbmH
dUTSs40tbsgMDPZG+EZ1hW6m5JXIKHBsOOiL/5c+wiywTBTRDHDgTPX4top883ki
NAzO3BZvK3C4tm9pQfeq9QqFrcIFK/M2BTLL+VWool3EJ3h35twYlhadtjE/mJM/
b39rpYsJz8qYMmVrgg2ODb5yGvH2HVSN7kDLmqeoGFXoa1pOT5qeUvhD7cOYu91D
pgNhHRLCagxh93yrhUK9lgdFRvucdFIRNNhGxnYA3lR19CT/oEJnPN3Gsb1AJPYz
XkKHxXvLSWzEUWdhh+f6XapE2KRrSMVgPZSbI9p+quKOIaUQQ3Ej2wBrg9J3+i7/
hvC+1vwjGakOLBKS/VTp+2oNVZQhPd37TwtiqF/+G5W48EES7N1IyJua96iG7Cqw
Rx0LwwLkHcIxwQaczJukt46296tBAowOVMC6FY+FfbkjDpxfsTcts5eUuvga14tV
J/BzRHjwqNJhL3iSH45Vpu6K8aCIPck5DFP0kO1dqOGGUZe0pPel8Q3Uli6tsX2h
UFzsfxLyCvK/8mXMugqgPkR0z4A0dcXXqBGouYN2DKNFIRM2+HvdkZXjh+MvgsFc
jlg821bt+IXqsFdQVA+Uqa3TF/GXU+Yrqmj1vLaU4O7glMbTgUjRRRWG77pjFj/0
paAWxBMnk0M8K6YERG9ngEg0W10xFf7YwGi19qckwLQHVS3+KbRLP+rMBfOLs8fc
Pd3sb9rdVnrbnihOvUmXKRpA/PFaimLpzdPqQOAblsu4lOuRoMqazU82NXCwDG+9
BjCJiDcj+iK4knbSLUBoM0xJ/P9WGKpbEw3yloT2RAixC/433cwucXx5WR81gEcZ
aBHuS/LoCfXEEAaYX4EfBCiTed0PhAX25gYefSG6Qz5Z+leiMkQOyHxI2iF9Z3ND
o0QniiypopCy0QyVoOh6SwwwBxEAq7BVyB31eb5057e9mP1n4Uw4vND7DgRVuiTv
XuXP0qJ0f/d9u38HyIYbf/j7v92Ro6rt1fqXxYqHQbcOtVgDzpLl9DMeW9Ii2ACX
kyYXWh/CAzk6SzYq1hGMiR2PhEQ6l7TwgG50cz/VKiE8Z1RtBQEhNBafCYV2ZD8T
nIYPJFd3GH7ynaJVj2YfjAlOe7EfWurfi6i2YjDfJzt2aix4ppvIkz/KoppzHyo4
74kJZ3cLQT78cxu29NNbdZxI+4kK0tR/VdBqYaEn1so/DDcpDun8wyPkLPsUeYcr
B4b4gRUOUbLqFf4PYWJoWnhuCuXWr4DVfxYtJOBP8Dghj6Q2MBYGy9t237yDuYnf
PVrPJugajEAWgloZYgKTnXLqN0PbdN279ftJLq+J3Xh1IDzJ6mv+82JXdQq60YxR
RY3t9mdNhfz54gQ0eR7MmnYBnmL8RSgXTuELp0+4H+7ih+Wn6RSGRBccBFU+8uvl
C4DdAgdMxgQTy2NFbbIGCE8rd0w0WIZQETUAL1Zk1al6ntVNvSpeNoUPbow8UGi6
NjkxOdjGfYeMBNQtwpdvUEE237hoXeW0+F97gEjsur+w1fjkNFVsrdYUOkoHKfwb
jK3AMTnZ2sT4ij1rxpyH+WCtS5kK2gg5NJZ5gphIKg4TXszehk+PSl9Krp0jX4E/
/2o7EUb0kKuRFnOsb7Gr/2+HwVJfR+laLUT8rrcb4CsVeGJH1LBObeNqk02mua//
DoxUQLejW+EHS9gsfhHpyGB/eXf7uc1SwuMAm83atnUH/zb97AgpNH2J2OHmxG2O
MJ0qi/0Wi8E59c5284OU+wV17MgOrCb/KIVc/FZA5Ng4WzoyuPrtoUHHeYzjIt2h
MmkHjcqomjILHDZeoRYZY5Y5Dq1exhy1LjYagwZMn8yJeJyJVTPM0lxji6LIYCcO
ZNF3hUhzdA7NUGJ3API6wdPYvOv0riaIwUg/zCOYVoAu5xkAYHznAVs47uVz32S6
i77OJV0ZclDVJCQIbGfIWnKd42+DuF3JLF6OR57m/7wtBClCudMK42Mx+yvQ2AJu
nlfLzqbgt36CiFiMt1du610UsV4RuI6SMWS1Cm9lve7Fo8Y8KG/8YuFXVcN0jRG2
7MMhGMQNgtlbc7l2v1Hw6Umc0QnqwbsByg6bwIsB0DmroSCC3t9bx2e9VSu9T3rY
HZVCk1+0qa3Wtm00EhCqp/h7iW5pRJDUfrnOVJCb3UkU0wsx+adtJyMxIYe3lhLZ
jqYcK0mTlJJn9w1/ctWNFYb3OzRyWcPC1tjYqsR0OqKqLCw7qzF0dMSAqnhpK2l8
bwVSMcX/PALvyD47lihb8X5teuvguTELaL5ADrDSOZ00ag180py3wDeMJ+rH0xSH
/Om6XuDBr1aLqMBaxGn7/jnfnGw1d9yszLKZonXSx+ZE0+yInkzKJFLjPAQAze2W
sMu/DYB3Z6L/AyxYoxQAP4YwBqaVDyQr4p/HC0pVX/h8GfRlqMIqb+mzZ/kbyw4A
rLRd2HbMCL0CZDWj1/tLpWKtcsshsmXJCimxCYJhGef8X8GYNCo/UoBpcwfPyNdf
6OoaeB+3WjnmycjH6Q8TGSMpVfj+omLAsuWUfih5j+oGbERZe+EZskOt3fsXwK/P
OGvjOJTr8jjNILiUw5dyutQCBSg/0k/Z2Cmu/CNkJmLWltNzwYKH3PfDYoPu1x18
m38z45oAxFYS+U6nu7ffXdV+dewfVRMMnGVeHs3sEgSuNutHa3vhK0sH9ODB5eXE
gN8Q69salltc4PYcAnm2BuThzJQd9z2RSGfDMLgaAadtbDAwgohX/sRjHR1Ek3Bb
suRZPuQHvRmfdTp+krMPOifuAVkzArk76qZAcYMB2mQGhqT46y09/DrebWR+Q7Xb
WJRfurYtbzcaqym55MExSE+yvPq9MjNgWmcIGnNJatJL7a8wLtnBOYToixXm5LHf
pGDZbEyUkPj/p7snBvEsmsLsmyjVdJkcAcTWsLzK5W+hDwVUsOyv3l+snObKec0s
AcvXxzjDSc3GymtK+7RZ+WWkwSDKTu4TOm1b9Gx5k2eb4v3kTAWMAN5P/kldya7Z
sqi9EUaNJAzLCp/RCgSEsh34FlujC8/xnWVihyMs+Z9vza05NWUl1RbW8IHJfUiR
GGO2UkDtjIfsV8EbLvLvO7JpmMslmEvDn9jvAQSkZAYL63mnHrJ5BZSBIsw0cC5L
zjzd94iko0RZPDPULslRZv+FTqvLs9r3poseTbh51OzD8ivQW4AI2QzU5ihONa0T
/iwIcXsuT1a3DSiTck2Bb5MF/xqhCW8T8fMvc+81blQAw7f0cQbrKsQPUlP+9aoy
tOE00R9htcic357OerTTk8JCGMboXDRirhmagCAjzUdvYQqJ9omseOBELgbo7Hzr
j2gc1ledFBxb3XpZXAeXv6wVDpccZjiA0MWV+AIv7eaBoDtU/XHIIiHbSY4w+tcW
H2XKf2mB4c6tWNvxWbe5hdB63RRhpncLEc6RLxNdM79xj3EmqMb2iQlns5GO9R5z
OgLwnaNT2SwUKSkV9V7wGvX11x5VJOFalrOJxTlG5Il5LB7VsmFkcShdJwI3aefi
Tetlcox+9pttzJoZWbwQ4kV64xCNAaRAv0gW4bgkGzPJ/n2qCk7WVYlAYtCjmYO6
jJ7GdDmm3Mq85MFSNmMVLYcLbdTmk4esSF8EMa/F8GvnbUbO4daiYYQhR1WJyFfV
omQyt1Crqye5CfWrHwDjbrIb2mHhxdMBvZfygGB4+OgCbd3DcuaTjK3/mNmOMy6n
GaBDjWJMt+VsWFhRpART1XW6geIuErHfyl4b4R+DXI3NpQnJYcKu+BtGKpTwGoeV
8gxSnPkyvyGOYJ3oP2xiz6wQq0wH04lFWj5EL5/pmR2qA0mKR9UpNP4orJNtjoiB
4Ir4DrbWIDSoyIhpTf70YzdpmRKNoHDK+lf/MS9IjCTSASDRF/17b/Jjymr84iZX
ApESPlEA9yjE7kCCf+SRMmmucp6m+ulQRF4VyuhqhUxMoG9BIKs0oeboGY6LhW4n
5vnErK2u84+2yKU11TYetVAbZ5jwmqvaaHz4ckiKVg6uYB5XHJN5OwPBmFx1M+1y
8k8aKlCcbfac5QmzSiUK7GTIzH1Q0dlgAWSx6y60cAwrtqNVGA4Z7pW+N+rftP9w
9hptXxaIJQ72Yb9Vt4eI+LNRiMiaZCLyN8HfgURtUbX4T8hANPy32BMsxNj7EFJT
cQkDEW3KPg99X1NfuBCJi4SZYAqaLwfHrqVaGXg2wkXtkz9yaaNjKbYM/NkFkAzk
fEsllTalFmeAqEwMVxArgOKIX/OYonCYyNbUSlgWxF0mL51XRSVWFHtuEt04KgNI
aM3/NLh//Pa/ZDgfycF6L7te78QT/uEZVLL16BKteTZ4MKZtZueRdjBwQvB0p2qj
J1KFWKK/7EtiL6GOgObVOfsNuHaRAcs1xQuRBIgUjlfY0wZZP39jrleReJLzwly0
c+eVhUcxXLMsnzVu4GGgfL9NALQRktqhHR0Vjj5BAqCi5OqQlzsfqOkcDcp6bYqf
MRmqT/QYLDKKweIs3NNl90RrxzBXFJQvQCYvH6dfd0SbZiWuhNslbEqyV1VNzd82
dmdjpv1pBOoHg6tR6vmbBl7LnnJgDCftLd6YPzWcRBKZj6g8RROe47saX9GTYvlp
hI6uoepE8sCQALZ3RXGPcLCDypnu0vfcoTq1YL9S97UyMOcZqY4XwtNK+XXWlxF6
xom0fo3ls4PdbKWNbw/ouOwaI1LCkOoN25cxW6JCwVmqm+XNwrbFNfk2O7i0VBdF
pLzXWhQfh0PFQaURJCZhhHLf92ukObfQk/pCV8v8p3Um79AqIlxs3kyto7A03dDy
qMQGsVMDOLjPfkiZPi4mbG7cUb4uB1Zt2/DmT8/NQyNdcMga95btAfX/8BiO0f6n
azTxtGHyjHc/kVBTdontY47AAujmXOYL7rPZvCnmWUpZmWQpn7KB8W5myEBOBOpA
PX6MqjRntcazdl0NzX277VPthumCUHyfVMseKokSDtEwVKnJICZsKW3MOrOjAlym
SxseiNDg0YobF9z3hVjxixQ/NSajiB5taVna8fMIrkkt2u359gwEfd4aSERXG3CM
Bn8D/lB+PPU3G+LM5LCVltxDUWqGdCY2p9wfNuqpx9sHsXtCwiVekGYc5wceuz0y
M28xZgSQymBKGpOrjxG7/rFVjhoIyzUDdnkHOgpGimfQjEPeNCuTN8ov6fP+OWYh
sdq9q8Zr+ta0HZeUfx0zWZncMHtx5MtH9Wtc28MYsWHzEiz5fbGFxbZO5gRpgMQH
DQDCEARLiA8bnUb7H4vgf5oE5f5bGW5rUMuyrK2lUzc=
`protect END_PROTECTED
