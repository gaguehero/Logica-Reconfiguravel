library verilog;
use verilog.vl_types.all;
entity BCD_7Seg_vlg_vec_tst is
end BCD_7Seg_vlg_vec_tst;
