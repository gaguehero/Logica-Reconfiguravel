`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbJeHcXQrNhMlwkJ1r70ND4FsEyRRg40RcM2EVHRFfUUopbHi9zkGJmRJAkKXHNq
AvhnZgZHSsz/wVUa1XHdoChH75JASl6uQlncGVpBCZdERiqsysO4vgRrthOFhv67
fTs7cRuKBPkfocwSRblBEj7dJeYo38ooARHNLVemDn9vO8rEqYUHG5xr5ytW/Yga
5mAKPfc6PFNr38HeTPmzZ3cjdWWadS0JYR2FDPWzExotP1F7cixC57CWFXbniIi+
o8lU+5mPZDRUJ3eHzR4vRAqUBSYDczUisaLiYMR0Bu11ESfk/dwkauoXxwAEJgMO
aSairbhgEPTjd0sS/ZHbNDT3chToFdvC5QCwixeopTFfGs1F9ZaxjMlgA7c4DtRu
7jXBwgZIyyhRQm/3Dqo/71YgjEyDYshqhacQWUza+ld5EznHZ0d+QXrz1tMYjA4Y
/1TqR3c4Y8LdpMQJZxEMJ1D7RBGpGYkysMtv8m29shVSCdE2zoBrzRJEhPDN2cSW
HpjV9J5BaB9v6avQctxbyxKB7Ij25/BiCjp23fIGmyga10JzaNWI13bpCEYUG35Z
bkFYlMPsMsjAVuYw5TsvM0nfHv/7AzzQdfAgXeb31RAy5EglXWbrTGyYslhF5tOo
RFSqQ0u+umh25WNKVM9hrRN1J075jf/dL93A60mN5VlEkIiAw+8I1sSBe7N3SOkQ
glX8T+oxReGUNMwMgT11dQsZryuixShk+EjSXUndVOPNcrQ4l2JoGubvHmDKHaTP
/sUnIoDtwhUKr0jd5IUjyQ9Lw0hxYiVpfb2oudU4L3gNARHKRq2kvhFA8Y0D2zFg
DE8QsKy60EzM0ET58mTWJ/TSsmbmTegpDxbppKkiVprzb+yEEdxJBs1pMUNe81Cj
MjCtYzkhBxQHRkvKovXZcxCRjFONq1/3RN+j/5yJrbEoiHDd2gfPjYsz+XhyjQGN
eXCi4y+lY2PKra0wQRtV1P+5GUlCSMjL1lvUtO4b3EGjAi6x0hfpCXDUWR8q/f/p
eiSIqgQyNbU6om4ftK5JT0Q5hynSOVOchkGPMLiwkQsCgxZAg8i7qO+ury8E30Zq
LZ6L1vaA2vCN45xspywbPQ5Hs9ORGlEAPZG0N57MxzemgSmqwdxaWSz1C7tbbKYO
6dpU7SWeGgA/aQ7Q15C4oPhr1jq7BGyn1grULZnZBG7oWC+tQ9BNqQNWg7ZqL23L
H9OZ9m6zDRCTx66l+d40KrQNOxZqqWiIQKZ0EdRtzKebTjZQ1x//YUIXJ2G9POXh
InY/VTFuZJ6Wh810azKa0KtII1r57zWQnftd/Z0Nzd4ng6JGnt2skZbu04UMf+Qf
1jVjNqhFqEoXsYd07kPodxAMTCQGKQT6hwPD6RdxcA6w4OtyJye/ag1TbJX7Jzz5
LTzpyP3BvABpnfT6Y384ttOYbk4NRi5ODLlOmnYIrtotVUEMLcbAOAm8g/D2ebn9
rZ1MrTgvLEh6YdPr0wx1t7BIuB9Ze4ol2xGG7c3CxGLSO0lZJp+8LwYlhsNypV72
9DaVvLAN1ipoUj8Co0Jl3AmNjKxkx6pNICtHLnndCEKGPwPlefZ0GitMwfGcQmS6
gC6V4nuiPRyjDkCgon+V+9aohEiVxxsvb3z3wGQhKL7lWsSYjV2vPBP5mdngGRPY
JX/coe6F+0Fu3xsIn/uHRCI8t9fL2l/aPFsAESQ01mt+mmw5O1yWU54ipQ6LK9TG
Q4ih9tQB+r8YHq+0meFyVxJ6ceuGI6E6sCneZVsIdTNRjr83/O8tg9L841d0uOP2
J6JVtI7yl8JWFl+E7ES+n3yihAqUoXll/rJ42/UMrpQJI2rWgLFTkqgZRhkpB2bP
0aIbKGyVWqzKfirrWKibL1+HsUF5z9eg2lf4gaFYmEKawhKYGO3DfZMoXZT2PaHb
TfLv2/oB99VoxYHIxQ0z2fceUtGc+hlF43EKLytUfXUZX+SoGtSHkraZNeTTMJzn
uUvo9Yhsa+7q4hblGQfI/QrqeY/XPWAlfAExlz1dVprbOzPC5oUDhufiHVe6Ahd3
KUDwE84p4QOZ704hzQKdwPxwfZDPYAOQn8EM92Kz5svAQW8GAK5dUXbRwMsnMwj+
vNsKzfm3VFYD9I4Uu6ntW/lT9CIJdBt8BJK+1KyfmcBGJECxlPhpgD8Lys3X5Fu6
LnhxOzT2xpFQC4sxpgq0YDpzrj4jojKHkXz2QDbnYEJ/jT6Pxaqac5y7qvKvBTCJ
Qn4mvLc2MOCpUyxzw+evr/xqw3VAjcrTlG3DZoKH8PjhHAn8LoAoGliq82JBc20J
HDDPgSw5zpctDnoOXvGxxIcPW8ma7nKEfWs53B1MpSp1Ghtob6Q5IjEioGvZqUdy
OGVbC8w49HJcLnIl5J8QAoudoqS9bTqipGTlj8bhXUxa0fs67EV/11HWWAietA1C
DAii4jKh7WtYwKqK4+ekOCOFRglpHkBE7lWvV2zMwKubE8ksN4KHc3Nklhy8Av3W
jkDKo5mcewUGQI1roKG58KT7G1NSbCIXnA/I2XMsa5VC4H51qK5gpj/gyUX7hhUw
D8iopvADb2Na2RbPMo0xZY7O6Vzn8mVzSccylcDlMp774jDCVSUZ1XOf5Fci79Ft
AAaisHyv+xfbHcruK5BdTdCnbCpOsRGVd7t75BBJ6lTOPCkFYxoUIjL8kn0crgDV
3mDds0fQ2scN1F2XM81pVd/czGYyhtlm9LuEl3+cgCdcT62KvvRUv/1HjdNkr/1i
P1BcV+EDOCAL7T0WNU+pP31WnBnmJF4qPHXS/7vtLvn/RAq+toF9rs2igHdoiOm6
kN/sopULD9s7Ecy0uI+LBLKrVrOEx42k9DHI4Yhy7c6IlGKnjBdoOaVG5UBJdlp/
Q9ODBfCt2Af397vKed482R5DJh+araQ5rSqRKiCCBQNLrOFwuWFjcL9j4PVhyLQc
3szhdabe5+++aQ3Ni5sufgwgKGXclehPWsMk0yn2vCCvurSFt+4JeBCdDAg+2Npn
UAbC93szn7xSHgpZofAYeHw+3rpdXVcGN/+EtAVtCfS6SpnT1s4Y/2zxAf7j4nW+
XXYmNwlq6SjdyjRRX/FWh+r0C0H9CEjBVmn1Ivimt4qYExyBABtBy9SjyVvrQ4Df
K73BoNQ1O4ortICVDPe24llTQovNxm5GQGgL3xftHJM8h4C/dPSHVPsY8nCXSakO
d4DnjJOo8ETDxFukKJ0NuDlvH+T9BzMxs0e62aAr5jK17s9AcYiNh/5ZoTxx1+lD
WHRrhmah+7tVEOhYVb46e7486zAb48JC3LbTK22MGdxh0KY4vLn2s0APge7KP6l9
m+BTw3ZgJA0HhRiCYUyHGJ1sFnbtR1NN3KMfddOZUqPE26us/O6iP40D2MJyr/M2
oio7A8S7iQhwYNLiXkUKfnNbnjQyNqOv28ImxYrAKeSBYyzPnpSvN0pkkKZCJpwC
Wtll9V7qynCICpu+ahvgINRHb40uWct+vvzbzVSoo3k/4UaUrVBps3T57fgwiuoD
1XHFj0WlXNotvGs+EHCw2Q7k/7XyzKq3jkxxZVES5X20JZ7e4j4FjiLF2IzNhAzK
WtwlQD2ZzDNeR5d0Rn87E40Gg522WfIzmp/JBxtpgGb4+nBds0p79MZ32G5YoP5M
gTJg+5cjk5wXfr5tJGZE2TbrNGo3l0Cva9wHDQlGEEoePkoLMvOa+e+y1B9sX9Q8
df/l3f2bfbp6CrBu624Hu6Yi1iggkYsRpuC4wA4d9EMeh6q2xTPXou0jZ8F/GpaW
/N7sqTXxaVVsizKzOYPJtIohKwJ4E2LLrKdH/AuAhBkRjxI8KNnh0yMfC8Zx1EXx
1N6Mpd3WjkVJxnzJJvkwy3qlZPCVLJA7ii0Gja316ZzvvvYo7vOMv0JnA8ALmpMQ
XjrEHCOYJjtMCmeXeo19vCo3Yqbn85oSQNUUTkUbcP6u67WYiqqlgFnuYhWPT/4t
ZF4xnUZEHf5t4yjTVdkyfu7CwYEW7GwfMlow9HaLneI64BUpmkuH0FY0OjLH4fI9
LJnXTfwNtctFND4GKfYSW4lS9cAmO5plYo0LwR+nz9LqjYqmRMpj69IOdwxtq9Z2
ZepO59BYQX8nBzTNF0hqySFCc+C1M6S9qSxbfn5wJ0tEyZZzBbfcVhx9p+OUrMIb
xqW9SnhZ2ehxDaD5l+9cp6+B0C2Wiw6xc3D0i3FG7NLPpa4R2ZOPcdu8fMjUcxfw
rIfg9zFKfe3c8t3gSk5nw9XvTAVGnTSzoiPQBUSFqY4R+opUfqYx32kvkCRU6hle
Oupgh61go+UsnbXqGKNYCQWin0EdG+f8qKatGbht9fVSZIHDdY4zbTNELiyxcox+
nOxASHQ/3QmolXZ2DoDy3A8HeHTKZVXt3nrDWXMORXWL7LEx4KRsXEjq/j0LG3Lf
+GTruZ2HVnBLJPRKCFBPUaEyC1CVltlK9BIb5asITnSUU2MM5mohFTGN3ld+ePX5
cbeGZ9kK0FDj53aCLd3JLxKHfnw/0t1nMz8FB7MPSP3od2yg+MaoBCGPQtIQGphQ
dfmbJkGStEah1HtwtaFlAajvmcSipRfAdtwMKObMalRnOnIkqRQwxK+O+4TEsUQE
t8g2ebXOlKS6XYQzE9ioqTYN/zVscMaDotN2Pfno7IwOKpM5YP0GwJJmHSfvvvEu
fNLcGmB+tELhTAlJa8i2+fwhxQdcnxvyzVRluRq+IktFSD9/BCnqbirQV/Q9Oc1Q
JKrWNdsQ8eNURF3OmWQjgB681Nb8srQKF+Nvpj80L9mCSCWnOeJib8zpxVzAFzBd
MiQUDjng/XlG9xmysW7plhmLyU7LmH2kYmN23ShrADiWvC6MAitcZY2txorm43Q1
SjX/4lfIR8PbTOzDjVkuu+xpUphbZMAQsBruIV++7AjPgj3MZgS2hOTJ3JxfwH8O
+Lve2fFmmkrDr2lgeJDorGPZ6AxAUcTqLpXisX3fwnMGdpAuWU6Q478aIOz/ewff
fQfiDg9YIjfExOS8W+BOsbn6/Afes2meSFnwtqCtDUqEMj1nHKH5F+Bl+SqkJmNw
8sOWvlaQrPH4BJPHAvkUi1DokKsGU28lQhRF4ZXUosC3ysr+78mlvqVp3dDBWqJF
mc4HNcU+LVIC0+GLNkcIIO4p/EzipBkElFEpnM9KZShdtzsr/LHnIOjDatkYBUtZ
LQkETAem8QxLsXZW+3HrR8EOCafyFUlbpxHthkSi2JLGWERhgGGbf65JL7ZeSZtn
pt616knWcbQIX+Skmi7gk24FjPGA4YDwhfeSN3I/ZxRHbah9wTfOh2pSGYHbN+6y
z5LIFRCS9r1VH8G1zd+r2kar4xxMjQnDrk3ou/rx7QjHoFcNOXTpCbCOU9oLnLQp
ofQ3kQjEzOeIQJcnxY3+4Bta6kwH0S+xWeUMn0zODyYZcau8pTy1nxBB9uEoWipw
f0kUL1u2eMnhBKFrP6oeXfjZVMAc3iP0gztWVokg7nZ7plksG7OzpPWJP1sICS6N
XeoNVGaOro/WNr1HEnAXLETz17nlnbbKOVOwdUDMpMjnI7ZkFEoXL+qu2Qn9CLDp
zOG/Xk9zwKo3bV+RFC293DqA26pMmI0/mAXyeudWunaGqP8O407fFKzuNIFnsdvJ
pFWPjoTk0Zs67ndRgJf9DmPrrelnFn6pmuibaT1VXdTKw5s7a9r5gDArGXmMJJ1u
FT48ej84gsBVH+KshCYVfoKOX2FW6snI1A6S/wwMcwSeUcHdRHo9xfYzmTfhw2KP
CAFwXdKHcd0EJzR17Wugm9YEahGyMs25CSziYKsEQQDE8LvDmYa9lLm4wUqczGli
P+Nppe8OpSvxWPqgWth4JjmJEhtaiyxc4Kkoo4hXL1PP1E5HSQ1ZAPfzRPSj06U6
QjidIUa1WiyLhg7FV04FwWGEcuNSvCm1lYEjh6INxLCH2TYtQ1XgNj1rPW9UAWtj
mTLfhUrStMFAFg0ryMO7V0zRD4XpBQY4T4dznSqY7Gz25JSOCTDZ4Rdw99hdQksa
Tcudlqtw9jnWDSmvqJpMquIOmphkxO11zT23Ju5axBRwcHKd8+NyG34QmiSOjHgl
gHJF2V+v7Hsp57KARZJKQxw6rf+Guronqx/02DorJR9hyAT73u6VJPE1zBGjzr8R
Nax8xRgwUNFWgvDgvS4ljp2Hh+4DM7k5o9y50v6p5oMevDYzOVNUtv0DHpHxFp/6
RC/uYdnlCBTe1/UOx2PF3mkTrnuOmm/CL7stHCFz3RwP/zQZ5kLLVer6uVOqvW6M
rcwI3CDI6FUeAtGCfHxGsQ5PoCNAlDVEW3LikkwdJIlfMoKIuI7Gi/u6dWMjwSG4
awOuPtNyjMvqhKEcwjn0n26LuFYAkm2GEFTYapk4UwNR4K62NIhP/RZCFb5HPZXY
s4K+ruUXI+kxAG9KS4xLZaJb5mrv58mpcXv/ruhb5Ong//Ki0ZrDKK5x+XxOYXmC
VRdsZqOVCiWjmxQB6nBQ/5fBXGIkPmhEdwDRFa6rlH5xrcUm9osS6+Mpd2HyBiW3
U79khBW4kpUEL8Hv/wFtDzrcZ4A8NwxjDv4qqMYAVVtj4y/fQ6xtj8BMCfe5y34o
xd9yzL0JxGu+Ze1Ghx8cdB63Dy4w0EgD/BoCabyu77O5QjKLj7xyT8mkAjOIisbc
hpf7j5xWk1eWtYmNm2rlVEVxI8XBF34kc+Z7b5gl4obc9U+hl4zQegQp3GhU8QwS
pKso9CmrgnsVIFb3KtEXFm+FZ19EPPX+6KCmcFQVO/YE58j55mSLkA8JaHGiDtiD
/DHmzIZ7nC/Nx/pazh8MrhIIZr1r4w9XoMb1YDgHoInM5U80pL1IAvW9n2fMhrJA
pagu97oYYlbDfe5+USiYYiHFAL/mn2azYNvcCfJlSdlG0zDiSqNOSil1HXGMGFzr
2PsG/CD2sCRd33nGB0U39gLYlUzEmYx2kgmRd/vfn6nVgLe1xeKFGGH25S7mAcsN
n1EbtsQYlLie0zLmnHC0qJc+Ia+j++yCxfkYIx+Egqvlc6L1TVsG10NmZ6ArNis5
HLr/b8d3WcXR71I7PQlKuqxQOs64cqhXl3JfZqr30LSTdswGMWkpmSqPA36RLGk6
tpPQFrTvNCQoYupkbdZ8CauyckQUuQzud+OMHn+Wbenfo3Lp7pJcnXq/TjxesFp0
pmbmQovkM6y4/KDjteppEFV/F5LxQVG1ryYyDm4rxQSO28ovorZlY4Hu4/yQqncJ
8RPcXZhOFGupglZ+j0I5ppHckZSwvMUjMwrzBzWSb/aSPia3v1FZgZF+7rs24/24
0cPpO2BO3tt4y3NIxpQLd+PpV6zX119mVlSNe6pCEI+PIM0xTTDeXVgr6S1xkliD
FXRwwEodrlAIW+yPfK1cnMI4lEJpFNaBRdBBOWnfPKV21Q60P4Zsch7iw+oSXhN5
Y5ySaYpRaP0iO5U3seGcS/oE5GcpNoAT/tN4dgOojWAiGlptbnHvZAfSzmnvvgHE
utFEof5dosjisNGP2sYvjezQOwygJUbn3lVHN7CmYGNnmU/FDRJhoS+/e8SXZaGC
EPjlw1l9B8nIr8JqwWZxYB3YMeDVGVWFOLcTrWeG/4skJMD76xejumkT5YTdz84v
gPmZtWZ7M7ZYc5ra+gAxdqScdpGIiyr5iWlNWusLbdgwmXksBYa/65We2wa4MAcU
/mQt4kGxn5lfgL2IUFoz3uOm+dQEhGpeju4vKO+OlwIfolg5DWx/k+gJY6gkbynd
zoqnxosfCDiUs+dcTaTgq1PpIoFXBZw4jgqM2Dx3qEydQ3gMxzZXCEL9oPBzrfzd
4jxQxxQ4UoflvaNP06kDrCUuHvvjqcCw7dmakK3ihTkX6Iui/vk84gricWYEivZf
r6LnyaaS5cwMlu+sKSKdLJzWxmxCDi7T8jE/LuNV3veOAZn4EQ5GKhBdYjGVg68p
PSP6RTaG3GM+0cQXVKCmoAvJK5f7VgF321ZSHf8YEjs4HC/T7rXB1Db6jQDktglD
9AlDTU0UB8kMIRVxYiig8ya4uDD7582mrfHVF+6XtOlC2gVDqkR+lYpHvjnehk9/
Spg1Hr1MnnYKWxzq6SlvKcekypCYNxL6diwtvGRbDnQVxZJRBEQBHe7PQfO5gs/7
8QomTWpvHpg7/vyrDkClthnaFkaeugZsmkAjVeQSYmSShDN5EVJ8bZFAK7cghgyg
r1UM8mcIUhkoE6VXHKzrsQZRHijnxCMQ6qhIiIAGXUVK1AHMgT9SGLysPkVJIppg
VaiyjPGG23UuLjfT2JYzjD3AEylDLG6ig8oJi2LsW2pWRgc6ySXCVTdQi/BtKTUx
fOswlERKqwapO2wqqMi/xCKqR32OSbto/D4jZYursWNU8StZVXy+pwRaBSXxZbzV
aLdh7fXCuHOQ13Iw2pHXJdWZDsvb9JJq394h5pITnz+57CKaOpkX/2gAqCoWJ4fx
jdplQ5e4TU423rILxwcSPC3CyuFMOYVMSIc88Ja3/Un1e4EkXRi4xgJSuV56fsmH
XdFQs5BF8ZWpfos3HwLQoIIWDbuClNNbHrmq/4p8bz9eENxAB6KWmylbrFnkKGvw
ZsHTtzJfUs303qj1rs/RCTTreU0gUHZL76ZyvZn62LDBrreQskkGR7kiSVyFC6Jm
shv/iNghfRh0UtjKPWZw4jCVAi316f3g0+02j90uwxev/IOpiE2QPK8ozflNHwYW
6preCbz9im1V/WJAEG/JM/1y+bAPsz0Dte8KFezn0cnacqzKF2kmv6yIeoPdifZQ
9M6fRj0dGDE1nvLUFtZKtIfd+xjkzm/yDbcD58w6LLrw0EE52b2qqF5bgx+h8LUN
CP9hw32cERghsMQFnnBsT/2uh+AzfD8vut/KeUv8mu/KFsvPTKezs+BUVvxPvHYB
XwZUp/7srn0wbdut5OGisx6qEf1Avrss0jV56YZbeXKoPqCruBVXIanW96cnMiMW
3ZyyY7CA97FH9TaurX5KrVHc/Qsv7a233NAzKrR2P5HdzmKHN+Vv3+I7BZFQu9ZY
gfSKFGIEroCvF8a4cepvIOb4E4/Vs5rfkRc94HH+eDstZk7zGL1Atqg/Oa/EzOnk
qyACLfbw8XTxMQSkrfLuMzRe1BtvAzZaDNLhNrDtRCOalFtJ60g73AaGLguBn+D7
i1ZpL9ub4JwRAgDJWnuaonBnX2RATzARDRGuaaDTgIz1ZDUXCDobdXQnUfcoCF7H
IajheNilREwij11Q9wC2HFZrzFScumBkoXfSG+ip2xQh8rE/m/oVvIYcBN70g608
r6fjMBgMIX00Txpy4EoPtgVJPXXaQ5rAOzEtogEf5tREdJn2Pg7L9xPa1zRwM0Uc
LJUyG8+GxO+GVN3Pcwtjo2WktUPi/OV3JGr/7zn5hPSv2QsvexVxGBq5p/P9sq3M
gpRFjeXc53tR0f/05MhGnBUXNfPiwRIdq+xlLmBNp7W1kjEonjki+px/ogNdKq2a
XalGKdY3gG6IxQ6S4x+GEdBXzaOMFjM2EmVY5Mj97mLCEmF0XPDAeJBRiCqKq3vO
rJf4ELSZzdMgFIw2Nl03gf7C6l7zk4Pqp2OZn8548Kd60/IPo2Adu55MKcQgSknx
Vsxuj8ymtjGdwD4DcN4ILCwC+tw9zjjxqOI7nuHJLhlTUtFWYK4lazj2O5ZCndiR
y9nRqJj1q1JBD9Tj8OK8VAaH8MOdMlfMEyx913/9RS2IgoZ5FCGAyRtZhZDMgWN5
NAwsNdD1p5KKW81Hed4DNBv/D2KQqaVYS3MUh3s6yaC4X/8f7LkzvpPnIZAWmprW
M5a0aKQvexSzOLL7SJ9h36NcHGQFUQR95hwr+o2dWwUSw59Q/9mUg52LuuENyXFq
7+FoKybOy3l+1DpPqsf/49QHPliwCWWtrYAqAAEE19p+tGVQUhftIh2u5/78Y2Lk
kMkeCBRfdoAXjGcZF4B9zJujlBZ3TSr7fWLSNzbg7E6xsPvV90UxpPApjjfx+KLb
rkGFYIj4++pbiazv/+n/bAapH9crp3Vmg/p3363CkAAVNUkGWO1yL1O0rNQAvWz0
E9GsuP5v5Swil5nEi4F0EMOYXhkmGgptgCG613cmYD+ZH18s5Loy4ewtuTdkWYUN
cpbrtH8+myMHmtiwTjSy10bJsCNM9vJSRH37wlrtKtEIDba3pV7UJi+6GKuze77/
EFn0nO8iRWZUpJbwIOOMhkAdY2D86dUTvJwXRLHPbmWOI9IL8hFARYuYia/TD3BF
zFoeHS11o6VCCWV04GRqFz3CVwu/yiE8YQ8kX3H1zH/8hefsRloC5miNUzcWXZAw
YcMhfrLkZCY/wCNYyTHeY3C9B8JpxO0F+S/8fkUWJ6DPcItftY3edEds0VDAjYca
PVFtLcWr8ozD+7r+0Ub7J9iD4iKbQDxQT6EGg6N79wQhW8+dZ+t4pP/p23t6YIe8
lQpOKLiAVA+CFqN+1F5hjOLad/AMylpAafo/gVXxiZM=
`protect END_PROTECTED
