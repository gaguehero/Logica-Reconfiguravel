`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8LxCdnVUXh8T/nO9EU7S2l2E7LT5fv9Nhj125VEL8ihdlW2QerXDwjRQXI3fmXz
7C4NCLP79T58NgpZj8RObemfbX8pinPVlfzTBD9F9lMBqGCgXcFV44tKS27ZY/po
mQxc+8fw0t+sskCDZBihNc9iMRu2QjNy6heEamaOvmby+nhWfuqiNqtJNhcGhRHP
RwnIpIOIisw9faunZjnjGk6a6aLcdXrFNUmzEK+rdRXYYKrKy8hGAqfXsOIYQylp
B7LU6Zza9011VnLKEl1Xa/YkJUgzSq0od6iSDH20rNlFIy07yA+hnm4o8kZDJfHf
A5sDZCiyVNzvEY0mQKGXf4WdjsmYUqnIvCg2UVF6jBontbv/NBV+RAfDfxJnk5Q0
htq92BnrGOOQWHNVbCHMEGGMCJuDQP0hAVqX1/hBybydo0anC3vQSo/B2OXY2miy
ryCnhDXoeAGnT3pky8vpa5echrAlYj+GRCCwiUXpbiB9DbuIoMT4/bQM4+WSxpsi
Cr/KHDg9P7osJXp1Lt3RYCgKEg6OQoAOqdrYM7HbeoZsrOCLxSlx3w6Ti5PTmC+Q
guoTD9LgXN47lfa60UNuh+V53BvnDJwXjYs/hxbCsAlFgNPCwfjHeMy0WUUOSSbg
S6Ztav4yK5+ByXPTk0kNwh0vVvYTVXEFfehUAbbokmoaU+WXRRKcTRji975TwHR3
aOGaH4fxdQEZbR98e+7wMaBBQsmMvQYs9NvWyUyTKuNxSLX0V6Kqxt2pGOU3XiD/
U1YwZynEMaBLHq844mnOQfYUj9UcgDam8/cR+Bvx6JejliXBzy4Y0aFsL4lFaXWw
ddlj6vtoLRn5ViYyMmP02jBWXF/01WU8ZGcjnAvs5Ob/dHkwiMBgfCHcw6gCTitv
bylzTuY46CZTvZ3uDljg5+3eIFjdZlqA4Lq+wjWssYY23N+W6NgucX3R9yw2ehvq
6s7CPpYCsBc+GZRlFeniVrU2jP4D446bYDGCdanj4M6uFukka3Sdov4YRtj9FvPB
KANu+HQjVTxAm+YySn5UY2GxTZLFQjCsgYdZH8SGvAyyuMuKNb4FQKuuKLmN/X+B
p78oKqDED5ZCKT373TSC9/zxMe35gmufTWqhzLP+j62Y0wBfuJdE2SJ/je7ipO0U
nm5ep124Jw2itydVcB9OjQrCqGXQcyZ3lJlqxcXdar5E0jZY6Pc6Gi5Qjik3cITy
ha+E4GQnX6PL9tqEZMgW2tcjYp22r6Yc1RLpxsPNGMTENzS3RORVZTn8Pl/MyoG+
8fjUniIx5LFNgSaGFnIeDxsc7JhP/S4rb59dyeDLCy/657r7dXGpuGndN6SD2wBA
ll2xKh33acMON/wGNMfsWNqKgH8P56BKX+Su5LDWNdMw1hgDuSV4b/3lzFa8uXbv
Sm+PiLDHNJGhlZPj+Xgh6To26TMzBRoJX0VhqW37ZvXI+OTsY/Hc0Za0zcVpbdsL
6R0qOj6djwBKHBRAXRysaL+PJR0UqPg31s0dGY1NY46A9gFkwm8Os7ZLipMUvljU
Pzo9DRrHzfGyPsKTtYK+17d68dPqwthmZ9jBrYlLUjOvKD4UAdTb8dDs+JLMNlfo
+69ILSQtDcBbfNlGV7IjeEmWBrzZ7f7wP3YLrLtB0OOGtmLUwlWSQdKvf6b1VABV
TeTv9sEmXvC8QI92Y+8gw2+Ufl26CD/SoB/wty+Ckd0r4pdR7o3zDz6plqABq3S4
KEvLrf+O2w6CdXmSj7Q1IxsyLDOkd6G+so+MXFmLCHvrKwMwUTkelvBa6WNmfvaL
ORKFnYHTdLENzTdfypZ+KN9xRRqoeW6duoTF5WoATBBcJ9mcmjhqsRzSrfI351sP
Q+VURJXUjjF/BwOEGV7ER8KXdD0kJXPCFtuwOgUyCB7c7DWb3Ygi79/LHb2CdUCO
t5je84KGV4E+9ogjwCQ5wg15ccwVaBQD2pdVjCL5rAGKZ5MDOKBkPyir3hxfWRfw
4SRyxe9azke5/2IymUvMo5JE6wjFC0xMYK47zsznGfV3JVY4A89QEMO55iIyettK
2L89c2rY54mnuZVBh0iiHcOsnrBoAv74WJmqGzD6pbqVlYVbL204lVIBvFywWr0R
zPfddCE1J06lenryN/dNJuutYXYmEQbJJGwijAad7WSQFFNe9KO5ltR4CrqzKBV/
xGSfcdLynJ9ToYlQCRToa9B7XkESzBps8q53AJBXNlp7EqO/wphm3DJTdtB8rjnE
nmcEieqjFC3PqdvvmE9V5rD4OdRqiKWTfu78HXmtmVh4lBakcA1g31GL8AK4iFQx
8br3cm/MxqozS5AKjC0zpb2PLKqR9Kys2792ac0/9DyvkutcACrXxOjouq9LVtHB
8TK/crDkYYk/u/ZqbmTg2qW73/6n+ymccWuwgRvgszZK77qiZc7YozpgptmG1+bM
F24pvQCQt/+vSDLkPN8/k6HPdeCEH+1u0l7XdflOsmnVq3UZdV8u0yK4IpMQjghM
TqWM90FrpuVdW98Kg6HL3RW7Du3/TPOMsPyQOss+leZMxpYcNKtc+hp0VEyQWXXr
ZDiZ2meRZrVA3/3F/CVwWPO6a6xhcJaEjPMKmSFjHiPpc+U1+LzeLzjFhOhS5dll
oJSiG979pEhuaWL1e193dEMaDEqpPlFws1olt4HA+SRnx5+yW5ucY2f5TJhWaTdc
kxGgkwHJgf7WqAi9i9RyWzTyyJwvzakepplcKEZ9RoPiDBXV4bD7DfHdvzKDm8sg
mv8yErO42L+IAXxDxji21w24tobN+xh2liZdGjNoUmtY4cUXBtkP++DxgTvqUS+d
qIqqDR7fBQ7y/OxWW0z/DG1rZ5U28hY4lnDzK8YbN6x7sWh5zyikvr0l95e17OKE
q+lu3isANeC5mjIpylBaNiZ8Hr5VzBdAGSP+VmlLXUhRvXBAAscIm28lWy6Wqg7g
U4AZGDWSPMg6wX+gHr1YgUJwYr6a8PjQyxNKISi9TobO8k9idqH5sy2pXa96/2Fm
Dl9LrWWwSM3QHg7odT1suqiKLdr34BDdv3R3ZrJKNyK1Wf/XbVoSFHaJvtqW4yqh
0UaDS5vN99JREYgR+RWgGHg1EoKKYgEXThETmiAycouyDqHjbl5Vl1FUhKXLt3Gv
TQbONRNR2d0L7iwkNCxqHuUu/zrnBOP5JpUYAewsuYfkr6nP++78W/Shz92Pupg/
nFhUOpt8qcT6SQuz6Mf89KqvCUYpgH5fRMYCaeoBNv35IEMwVZgYxqlf7znBgdFi
X0x6e7y7aJSbQJldY31AORXKJ6kP+F3MMUG651ImKMWyxOtpd5NStv2VCDjHamzq
fVvE2h2gSB9KQnMeUxqlviHszwQpSF1i8N/f+IUJlK5Gwm1H8IKIhlM9k54w0pzn
jdYC2gY1InPGfcSNa7lu22zidy+YVWfBH/z2oWcKOJXFfTb5zLbk6418K5XBJMQf
rcQV9msH+evGdMDUqYhaEf/0IKQc6KRiJKJND7N9fRtZYDnZUSCiYD8nuqhr/evZ
vv6T5MfBgMKVUVzXATs1S4z/ZVemuIlaNtwzZCEOS1VbjrNglefq+2EUmlPumxeb
m5kVKee7RrvCQ7XOH7TzwAl5woAqu+AdXbIwMffZ4sl7uZMkphJduYiTz3goO1lj
zKQgHB0WtCJFY7qTFIYw0gE1c2oxaTIBcHrfSkAzUizD0Sb8hlmXOPeTSyhSQReB
yMNkuMUWGI6F8TmbyLMf4+KDPnxGcsQ/lzE2kndRH/WRzvnRQtdQpEbqvS5X500W
ssm2AAT5q18oXPt2nxV6AZhWsuvfLOJpPHGqO4nt88i81+o8QJeF5QkeWHwsAWNm
FLVW3du5/+Gnlu2qm4aXFnYyGYr+N7c/DpSymjZdkwn6CYhFfKA2q+uxgmXNSihi
QbXFGsRfl7VlnAKVe/3/bWSItmbf5pK9TC+jMgf/3dq94KN4rZ4XTZvx+a6zviIB
N4qTTdoBWaKkFPrwbcjIYy0LsEZ8vGs+ZpQOeDQQI2uVv3qNh1OpZoOHi1ydkr8E
hak+Y3nA+bZMGd0LbCp3yMN7itA5ulEO6Lxac4klFnfsmQDaVPhTDdM0HJISZs/m
4AKqik19LJZPfHtNsE9TEbFXCSfg0DOF1aaDm6f0PbuQ+Hgy3ub/QrnJWe8/OoAf
HkygR8tjyy5Aw74QYBFTEP3GFiSfmO1kkCBZSIQzvq2nkztOdnioYcnOXQ5xBAHs
ErgIZAXMmHVrzPDRjV6X2c/klQVIBJFZ/P5jJUbuYcXTK07ypfutr94n5Mu40Pd2
pWt5evxXwnytzPiJX2izlt8FLgMDbENgCwT3pJ03PbNqnGtk9LhQb9Yxpy50Ahxd
hKXL3j0nIvhYCHwAUVNobQbM5QbvHTtw0V/OW4JYnAzoYq9Y7Z/BFqbkboKdKVLA
QK2nbob9eX5fBdYYbla4AoSJeduf0pVsUYmPfrRq+m71TGs2vqmn+L2p3jWt5bKg
fcNhcpj0j95t7IUleDaBKK6C89W8+fxLz3y7uIBI4mSJyzKtQlTYXfA+vnuaGJp0
wBEb5V5fTAnJyq6Skx4fhY7ceRBOFPNtMZOGqblUc6jF3YSRFq36xgsdegsl+bMC
UcsBuubMCovc0BNRU9qUNtCK3LGsqsabhOynEmzwx/6VygK3AKKZEu7Texb31lLq
fxyRtdXkKnGVdRWeQGIWomvseG0Irwv23yNR+mdJaQzwwfayzOltMaAPORbIDsZJ
1PxTrZjimc69q6Ou5NE3ZzkafGlSQsHVTWYoU8/rNDIjN5dbnwHTgUvCnCZSOGXp
BjvzWJLmiZ5d9cO8MJpCdQNMv29gtu6qc7ruSgPq0O0ojDWbFyT9V6v/BM5CaaKC
54/Uh9OB7XWUipYc9VzKZylpE0dxo8sW16IujNQPj3S2bCiKBrjO0Q04SyR/GyOA
kWpGdSBAud8OEwcMpdHssqGtCvnmz9UaPREe2sicFfQydOchZC3VGUtXPyI+e0Co
jxF/3qv9UW4hbeDP0a2T9sCPhj9ePgkSwY6U8Fp/meHu4owuJsXlMZFQyyMcwOYo
UNUX4Pa1lvFhJ+zIF2E0Yyfd7KWRfnBiWPMQUAbz7as2v2QhyzmIyvvBqkgODRRh
mYIAvsv65W+HSS02jlezfzZUo+sztkyD8uDy0NJk6aTkU9tq/ZiWivB9tvnJuldN
OLj2aGcQ+ZGsSd7pBeYzVdEWn8vDmH8R+BxKdl7NXzEUyGzSSGdyIsIdMHeBP2PA
OG06EcKkxjbdYaQBudYXLSWyQ6yKn3eQKltX10DNKbTagNowBwhQYKy+la+JiusK
DPuAIv+3udgdhuKE+HeyAc6kEc7LK042GKIwSYpCXaFLtD9MWuODHk4k7yNMH1J9
W06D25fx5jZRdSYNaJ/VJzMPcM3EK/kSEO3c1n2K//zmImJl6p+W+tDu/uT2OU2B
MkJLEMVPbDdcUaHgJ8gDUafi2QgfvQvrEGPocGpkalWO75Nq6ajMGkWJL5lSAbC5
5CZsd8PDhNZGgSzVSBOcs5MvsRWQmG+gBOhB8aV8RHtT6dOokudGAicT2K7CtP2L
1ZuSmc2Zqb1zxLw3jIizRM3niE2P35ujrzCh6mmBuuCcO60BS+pjE6yVn5MgH8yu
YMJANLBhIwm0qh8aV83e8bcWQwGEUNqZmcnaVsLCl5UvQLWSkwjNGjcqz/Y9O1+o
qapfGWCAg89Q5jp52dWGz1W7jONqJobUDTJSmuO7DolzaSYkJbQ8koXycqZAWwXh
30pkbUVVpXowhAINgTHCnifuDTP4IhxGrgwriBrm0HHUau9G18YkPwzwhHNdfGYN
Y8lKnIgYFwKj7eGVxOZLCbdGhuiddpge2wvm75zjy3xoqH0S1rWJTObCCm4B68T7
Exr+wUp7Uc0Ru2AUKXkKiUGwup4S3ojk9sTK1vvYZm0FCkhzt+OX6sZ37C7uk/V2
OzokbBvjaUGgl6AiQ8T0LuEkp6JsO+8WNWYM3XrfUa5NTdx4rp3Q+UO/1g+sE26Q
RL2TwWGCOfZNz25wsSdd/YwkIEbwCQ1h4bTLdI7w/JS2GWXvs1ZsnL5pD0j0cJ2R
TLNhsF6caAXjV8CybWctMm/54HIhTN/DPTmZgHvo8Rgd1PC87BjRqJoQpbQFfMZ+
p5OzgmMUa+HufUz/E7QGad8wMssbm8gIbtBNLZU45hXzp0Yr0wdYqlkonMTpufTP
Tz1VjCdg+30lK7iMRtSMNhhANAZWPc6YebGfxOIXEYUnjLqXzZz8sxbpQauLo4e5
ZEL1xxk0cMg0cQkCjpGGoZrNWeGUyC3VOCTNLlRaRZP3HpHJWRa+S5JNln3HgUrx
yJkCdY9uMteHRjG4z0ftTKQJh43VJkeHgD1rlX3+Z04Ff2tDpqshgS9mdj7WI2RU
d9OVbzlIRONNTtTtj9I+DoX0LUC9HtOmPzyOkzowJqk5L66G5/xhmZa0gRB+rk82
KCU9mZ37uhdeTrc8znGoz/rLFsWv09JhOp6TOt8iatuHEZxcRedaxa8laWqZmOhh
zmhW8igKpfSfv74+bnQyqFp1TCV/sPt32GDTmW0DX4Zddkf2n8JNXfJzf0kkxf3d
GKllrD1j/HmkT9WTb1hPTqBp+SEaiC6G4rfEu8zuMJMEm3iqumYHlgWBdtgwRf0S
qNZjAAMs2XLxvM8tMBhDcGFKZj730t5/1O5DwsAvS7sMq+EV7Hdw+G08rEERTaiD
YzanPxFCBFv++jZHt+xC+WGCjVrNzNlQx0cDsDfPo/1LeUUPa+5AqdKtpmJ1f9Ao
zqX/3ZHYVqJdXH3mYXXVoJDmAsE2vdpBkWQQczErkZ8Ue47zSctNsT5A8SQnU5UU
e64ulIh7OQPG4lvo0Pp423uSvgyiGfiLOTSyWEdrhxtNwdSozfwJmeDhSor+fCTl
xtnEDuWprTVvCf7XvX2nupLHgYQvu+gHhgFU0gPoGqXAXiyEtPr0WXCl1GpYnGRk
2+8JMsnbg/6P4ASyBMldk/cdnw3uhIgoo6cAJ10F+kAaap8KuaSnwDF1ZckHvSII
V+NPup/55v2u4iv7xafTvLx1+KsXOBcQoePINnjhMerE+lrz0zfU9ezaikwGCWoZ
w8KZwfBo9p6gZDUVdYcJXVrPChFZBwdrpZpJQnKXYIRI3TjV7rD4MkJwJqS4IWoI
MlnM9ifDRc2jIhF0+b7LT82nDPPBlxXYHs3pkkFOwTwH/ip8jMAjc/WR7JZsbIVp
T6KSoIKEseJAe/WezjvMhbaJHwOKRjUZ+TcykJPw5Q7DEmy5TSFjaTnuYBdkQO4M
Z0LN190YGuDL70LBpA85nqUgX3qRWCKkB0XdLQiQJZOUijvwY26eBHZ+4SkE4HKf
YafrxYAIyqmoUv6ruWfzR67A3zDrTnOsvi/TFfhExU0ssadIxghiL0AYNZ89Z7yj
7kF3E1g7YJgnQ5Owk032qf1rw1P95efoaWeTYyBU6KC2jVqI/yX1jyGbc0Xs4PDr
fqFIiTdifJ0GD6TbovG9/9GHK1Dk0k7ofZdYmeH7fHkXKmEt/UqrMAXwd9aLo6u8
ZQCZfpTTpbcWv587qumNApUZrUDdPe6Z763Vq0/EdL9EBeyEDFf4pm516uBn5T/u
KDYfRX6TelS+UNO2WeeOcTL7yx8QkYC+IYlWqP5ZGbM4Q3HxnIbqzdxTCmI1+YPv
K64PXAJNIih0hm6djU+t/CPxO9UGNKA/MALkzyLMI2hIuqHCrW7ySeDhnrNZYrpl
DsfmgudTTVkVYXKnExgkGI6ckLGnqHK6dAM0YGvxc/8xS2d9Zzr2AXiJu2ak4ucd
DKyoUwKvA9DCzxoM3uV22tb+wEnhsBkWm1cnuCKJc+HR5z98Oo23D/gsX7dUJrWM
FX12rf7hT/8vd+VKz84hGezpB+3V7xoeYAe+k6GFXonLHqED7TzCNdvdn+t45pWW
DuFQbBC5BZfzR4EH6WYMDsy0dJQCKrGHAW+df9UGVXaSVKWWxX6ETO4KpVLRzKwF
HAyDv3tE1rE2IKZbSys8SdMScMjxJsDye5i0y9XyPUCHFxWncAf1H7xLtcfdO7ZB
bugLwNrP+Idq8SseKH/SWwH+K/aI1RJ9bdl6UMRlzJNhQGwCMBJbFd9lN+/1gM/5
y5uPbgUHt2MBx8tUNL3Z8uviYQtS2n6Nt5FtvZzbQXR5K6RQUxjnER5UvI3f0WcM
0zXVcwvrKENDX1QYDCAbtFQqlSgGYSjoxyDfIW6grg8/7JA+KsYBIeSvr5ptK8Eo
Fol28U+4Xzch9yzhPOR2cXYOJahga6XoyLIWX947vh6WtzJJ6vgoJg3eDwGZFaQC
mwJ+Fb2ZE7raszHhDSCHv3eew3QrdP01t5/KO/CEDGwXJEdR1F4GsfdDHpUITTH+
r656fUqO9MkXh/xKMhzsFtnln0sX+cyiQ33mYozl1kuydXcIuq7wFUEwKwJFNjA3
MJMSr+VuY9ad62iKufpO1p4Ph/RuvDnHP9upPapJeNCzYYvmKC79n01cNa+J0z9f
pgdMKOAx98XDnBr01vbNNwr6rm0vBSAS9ydsmofOay14+8rbapZsEEnBeZ2jnQ43
MZFeiKcR6H3vKTJadDvh3DNu3E194gITaxEQUPD63mhcPhR8rbJjqMTx9TiK/eOa
kAGnuoezt95tkhl18wFoO7FMXniazGv+jhthxspgT7HpxYnGj6C+16ErxiTM5Hog
Wuaa1tno9nMGI2oxc7Vp3coLYdQIOCs9nUvryVxdqXIrVSPBZ0045GBy9KN2pPf0
1ogH/u7RcDRsPDIRlslkUb1ZK7hFX4CXAbgL8DwMQGvrMZpAuu8WF738kjt1yK3u
Wocbhmr/g9COH82K+RVK7c4C+o3QDEDNLaN79MF5cuxjapKQBdYZ/sjcVnJ51jFN
oNl3/Rjoq+v5nzLfJ3D1vQNyC7D6AbuPvdqW4Tci+p3qS8rQZcX/T//0fDUyB3Rm
fVm+9ZUVU4e8eblFmP0Dw270pZAYF2viHM3zkWRmJCYcWXJe1h1STzsnMlPmfLa9
Me2q8NwQkyWAafYlMKJdILUQ7Y2n4G5ahaS6zpFkEPuRRKgkktu9VYIyy5MyWszv
A7RzmQxZfwIdeGQlo3a+eB00ljx0v0GqokNEX42wlmUt+C/udmI3k6uR/58mduuu
N6WGnoNIuRXWbtgzxikbazLO3kw5NH1QJSZYXmElPMngbofQYfY0SV5R7PxEPm5Z
Q5Asqk6tVndV4hC12adRW6Tf2r0aaKu5iF86C7NFcja2kCO+YKtj84cjsIypjP4t
3Vbgo+1RMbX8S/kL+A+u2l95mHn7O1ExztkF5n7SKbzHzcBBkaj8BmjsOIJJ4GVc
ZThauI2pTwzWkCAMVRz859wavpXJZvjogGwNoORLApAI4/iEtXAqG3tUt4SHDK3v
pPzCIDmA16ShrLVqSdrGfg6Wl7ESB8rUvzRIFJjIYYTf3ViIzI4iFlvtXAAsWPrY
CuGjSvBLh5KFfiXL/g5Z9L2LBm/XCN5x387ppKGJ+egzWjQhsqk3GlftbESl1ck4
wXTfjsKq0LsHyT6wsb3mjtXRAV/HV+rXuE9I9VjW5X18qLEnaUNfrfwScWn+QpRk
jDT/OoeI+Fka+FEFp15RsIdELZ04GcKLrsU9WVZXBjZ0rpuY1ErUOQBSMB6gBkT2
ipcHj1n5AoaClDXdKgSq145LWBBU/DV4sG2wetLDnvOkmFzRoQeA/rnvIc2qzmnT
EQ7asKFLm9EV+jORTKsiaNIqOv/NHS3Fh6a8Q2Ck/IHe/JrqUTnacFRpVwwGIcyh
9yQaiTWzexPyHM/VLtxjiGwv6/KrLmn4tQQH6EKSrEr5KFrnr0Cv2dEKjozIesIA
MoyiZ0v6FD9/Rq4yC2ETOZP0g80XAar4WyoEXzY1Ww5Yc/CuXwDCuzsSQyiSZm3S
kgecRrrmxTPF3eEnntpmD7pe+gYP3Kegxrki5e/vcK7C+3IPF8LnMcmJ7FAcAQU4
LrpraIdZ+JcImAlukCyZAZ3bqY5s7OX+4AiecoyzCwmczYC52tK+RZnpMqO2Khru
PWbqpHYxBERXdl88WvBSY0HdrP6YN+eVcY1X7ObfJd9Gmf/nJz9vRlpeEc3nv4tJ
YrQJgle8oVMDoIfu6SOigsC5HGfcc7OtRPsuaaLTt3QRpDhyNVmMqswXV5bRYYJS
s7kEUxPjeOmJSxcXeoQScAxDANnS2U5PK5zHpuP2DG/cXOY6e9T10wnCfnGLWPi4
bqZmqX4B5c2VOeUTpmcsfv2OhQhYl2PeDqdJz0Z16LjdaU2ySpz+fV8EY+vtYuaQ
gmRJeCAX9UJhk9NPMMpE31MiN/3EndIHZ8MsrkIhhe/WVgpQ7rhOj30UdXvtRxsB
FH8k33kmiOGEWR8vUr+LCNOju8RIdNA4QMNDqrHHsyW1+o6XCZA7UaeFW+EFQVG6
PwON9DA3OFJbaSRD/aGNs3NZyIlAbbLWeqH0R5GD8Oc=
`protect END_PROTECTED
