`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Hh3t7vjB8lGswxc7CfSZtEjtF0QoT+rHB9vzHy18ZR3QQb3khW6dgccIuELCmjK
T+65A7apMvzhdoPgSn3vVFGLyYqMmHattwmFETmzefNTMZDc4+837660+VHLK8su
PgPDdZXH1AJH83EW1K+R8QesSiFtTvlcTJD6IEWZzqOhmKRrGl+0WqtZ1IFspe+T
UUI2KGvwNGR8NP26cQR/f1SrRp5hRP1hehIX/JfwW1ccFC5AQS/3YhKv5qk3Vynp
s9VNs5KRz6fujDhFPHhv2Bam4GquIKkjI6nWDIi0gR0JYt3s1rGJXnotsa0NFzTv
87c1WLER+xLJ2xIH6MTZ1OE5+Vx19FEldEuhV9s8scvPjTuAJfGP3QYgUwSeDz/K
7Y778gagHa6QfZE58ChYFg77iSPAmWBw0OipahUivAF2wLI5e9rdBP2ITh4Hhp8M
V1/yhx440aJKvdqhHOkIWbQdO6EHw0aZL1hxeBwvcln5OuKcHxUGEuY77pePLVZT
hoZdRasQ1qCajNaP9Wo+nfbcItIfkVtPHtEO7X8WRnGAKYmIPiSAOxDtbp3fCc7P
GZrW4MCLgY05u+A2bQmRt+m/XiVhjb5/l2BogULZZsPk95u7+quKH0f7m32tZ7ju
odHG3ZZVfQpkQ0njukcZnYG8fNY9T5LuD6hNg7rSgWIlIMo7Xwo5bvLF50q4ehXX
`protect END_PROTECTED
