library verilog;
use verilog.vl_types.all;
entity totalS_vlg_vec_tst is
end totalS_vlg_vec_tst;
