`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCz7aHFubT4xnFc36aCtsA+etkc2EK1KPMt1BzKu8eoB4hxdqx4Z8+/LF0JknNbR
gR+sBbv3jurAzRiABiOLYMPXW+fvVuXnugjYaowK9gAQsDAO3fYcoJsB3g9nQJst
5YFPmEyY5qqxz9T57kKwDOwslksaKho6bCPW21swqZg8yWfVG5O+Tf8e1THNtXJ1
dCXfeBR4vISVnLAMZT7FDZEono+7Jn6QDrl4HbThDskVDdwkaLCRcQTFxgQYltZ/
wsZevZJHXB4Zu19ryn28pOikwr3zUBt956cMAFKoxvGoJA1Yw2Hd8gMejeaflM6n
jZio+/TX6DLXcZsJ6jiK73ye4jzistkCol2YxxtExH1q15JVr4W0EU5HVEdgPwdK
z9XTM814XP+jgGNoGDzfCCSFrvmGG/vS0LNwuZV69qdNihrbAPiO8NX25gHND0gb
PAw2ZnJ4C/A2Ucj/f3V+Hii8k96yyPoZx999JIK79DE0R+lUNQWkoY7mnds/nYET
yiA2LW0g/KEO91rcc8mPJjKOAP/mqIuV8bGH2Rz9CAlCIH2fodVohh9JaZ1kx68H
7QKmGWEQLh0A9WMYSrmhZbwsCceTZENyI37RAlFoVgFQxoXnloim7n1LaaQzRDCv
gfj+hZ50BHgWq3yHMtli0WKcFgM+aQjuKzN6KecD5Ul4qhGDGK/CL3I5VFENaR2e
kaxfpf1DNMAmfOWg6g2qzed2tpA+zxwF5mqXbQWPdQxW/bs/XW2ypT5ti5NiRYOe
BSaHOmdwR0xl3CqRLap9HE7KgF94uep3KXaa8aDF61ZBaX9gz6Dz7NhsVMWkEt55
lc85BjiSrpXeI5GWyUEL0pBIiKthgDrxFtwD7A69MRTK9QRPwZeyG+rvkQJMwO1n
2uLqsWhRynGSvzwOpCxpdfCG8YcTdY87oMYW9f1pqTqnJ8Q76HlTjUcLsJbILV6I
kmSCX4l4Sv2HSl08n5cojnKeI0CehhYdAN0QKSK9sTr9TNw1zc6r1lyTAxMG4rf1
KHPMca14qHaFDNLe3jMuEhL3IjeiQSuBP0SrQBZ9AyHQ+wdk8Pmx2zgBhLnG6bGg
VYEOTsMgSHQsh4lKMqf8/tbj7XAXRkGorlEK1Rzmj8UqgSeTuMiu5ldoRzEAZGQC
zWuCjRue3BNOm13MOjX3fAbvLrujAcXE6hnvZxavugL3mdA4gOfHk8KjvB6ocHDP
/XjqJJ4H5PZE+o1Iz66ULwkPyDcN+LvaCAoPfx/0QQbuX0Su3UMPn1yRluesnkZU
koC1AsT42lrk3k8i0nsFKDMU4OhV+MTsQL2CW9zG/nZNfiuUSClnWjtmUDWIqX0r
t9+gI8p2xwPMgLVn90CLDhJ+ZMYQtdb0YrfoUT7k2WMdSZvj+0lQcbwWVLBNIZ6y
yKzERzIxP2FAAq9m0AwHUQOqcPg5+4BwOC4DwNZaGyFmjtGyN5l3sMY1fHJpG3Xd
LcA4BDoDNDcv+y8P0Ar+uHY7qKqQhhqeF0pZwmsH9DWG5QC4D0IVehR/BXsenC0Q
p02CSC37D2fssghMoCg+lwOmfd7hLpvM4gbFrXbSqEaWhKNke4fa/UtEI4cMb5E5
ZORe+30CZAIf4M0zoTJFXu85s77o8GPJusZKZxA7HXK+w4ct4KzkJXnid4DCvJyX
RVcJsFAiR//5Yiam3cOxcpRjw4vAvxkrwT+r9eOpya8jtFkWrhwBnKmKLV+L/GYD
+tD8WMSoMF1V0UoshPORxAy7IedyfL/0A9XVEM9DE2PjX5poSZVvLvMd32w89hF1
rCVLvawa0KVvFa3lXCdKAcDTNwVXfJLEN4pgae6sGh1o2CYi4EMMyQTfgJDiefv5
OE+9QR1bfhe8i/kDEjXqyoR2fBvJBAuipHgb1qJkRJEYS08PYAm/AcVqD68TIc2y
0Jkq6aEQ8rHtKzUmAZ0GOPDEkhRhkMSWEB32oAj8auOKn5NlMLsuBSrW0geORTzU
uTkoQPq3zjWWge3vBOrSHSJ5Kzd+7pxMPplYS6NVIYXLxuq6+4Uf2hHNHjk0Ous9
MGv/zBHjpRT636qJaE84gD9N6InCc0pU/ojWsgtXHVes7R7N1pZS2EIQDalXrmNN
O2W4/TmMzvUpbosHdQMVkrr+NkA6a3yoEqUeHE4r2DrcYeJwTf0XAY6+5z1m9q8l
h4CTxjgW4YyG4jarxky7NiYzH2wS9xszEGXY44zpvp3PXvYleWhTCAY9yqyFOlBc
FXJIw653MF7sEgQVFL5Ftq/zN6eyp0AptuTyKaCYmeGa3ag4cF2vVmLTwm5xV/oK
60ZmoDrC/GqBZ4XnfaKze12yyRZ9UTARfIvvF8tuVSw+0ZRB1D9cnZMNmXDRhG30
+232em5KyTP91hXu6n7jO8WcEH+bpCKDdblQ/y0ums8DzLZyRkOVJsDI9PtaMdVl
mgA+aRGFhanBvlJp3D4xzUsPMOW9ub3dYAjABaIamvql/+PxK5KG8NjvGzzSwFea
Oj6IX1KGOaE1dyHfMjS6IHaK1p7dDIIW+DYLBkraQhwTearwoHY/BzVbGBbHWOvE
zlsVkUWitJGvkDhZP8owVCXNucLAh+kjyL6qcX2zlmYHtPm8JofjQ7Iy0vRFY30t
fykIdAx2Z5KIltMlXWjRG2N5ckFlJPAITxgBdKxnI8zGzupjUiFxQtJ3zCF6Jad8
IvV6ilO3vFb402QwwtejhVbdfig/5OIo4TqRIgNZ9Poi6PhPgk3Stp/VR/ri6k+9
SFBsARoEkZsiGcN3YMvpTFxRP7ctbwxHvrxqVRyKraSSMuGnWxtc/KE8eO2PewDp
eeGh6Co53kc+OKS0ThSeEBROrwKfACE2TH5d3IsFSIEUpdqVB+mzV2AfhWyXH8Cl
3MJkE5LRnons4eApG29rHQ2Sqw3HPqVY8+G3E1nYlt4P2+WNydrMFM6hg77KvNnQ
Jys7mIXaGrzZv3FpcxputBCP5DyYHC/ZsTR7SoLANjzvBObaS9vexTyD+p1wm5n/
nvnw5ynD8nMYByKCjrc2CgVVPZQ/UE1Z92VceIxWB9tjn6ZddPPpg3MiYyuSwthX
Y+5J6eSNNV4hlP82lbr2izXx1fV1dAR3qEMSr+3HY8IXCZ5TnvhbfrJKMmvuSr3s
fDT71wHgNsk9yESY17zxl1yydQd5py4x9JoKAZRJysC54tpM2cxfTwI8naHVYGF8
yWqgB51Xwdok1PrUb4KvAkMnp6j0PRYWYdZrs9lyAKuYsAILuP+8IPhWx2l6NR3t
oM895frwwhAIRxPtlA6Kzff+wc/7C0kC4wmhTzyScHtMmfcgrmMPnnF5sYne1zge
UgUkScgnbM68fFb8HQYH/M1cYZlbgkbYKuXuw8FPvLgPm6CjCqGE9ldnP3QlzfP4
j6zTB21eCUT28VjRI7ymqNukbQ8nizzcVkzu312nUVPWx5v0Mv58sJCdKR6v66eD
L1RIgKK1ej+5ormwmuod+Qw1Rmo9ewq/lo/DIsyBogYKD+exPu39B4obpT2mHtjx
NaxkAQvedFjo544rJbZWqCapmVjTEjTGUVmN0iJ+/9UleV6QSSw4Fpv+aBuUmLZ5
Izas5fsL1VflxyxGE8P19Oizs41bz2dOQAJHCqeClhrXA3yAygd/p5R7w1FwE8mD
d2d4LGST18s/7+5Drut6t7XbA0zmXIg18b3tEcUc3Zm1UqkaZwPZ+fDbSSmE34XU
hmD6BQUlfrwjZ4wKGUtZ3SlAYk4NjDm7aPaSOdQSZIK2zIfr5S5DFSXM1R0e5Yjk
2++rX5MvHk04einSJ3c9zCsK4y/ncpLt+zF6mJiiTbN16mp7mFogirvA/tjRyyjm
VV4h+PThc9ZI3FcU4fhTcQsLHjWTz4sOwPBjPTMl4ZAxXqOl+lg1gO1iHDfqwS1v
Bj7RcZT6gNfZT076a99uQrXnW2Sr5WdAVwjEc1Bj3GIbjUsIub17562r479baSxy
rC78aBy6oBYk0wIF+TlxVj6MLFtrPGN1OGtWwwmXo0ukfXIBnw00twaTKLxzASr2
46OxdP56WXmMSUXJp8OdaKbYdeWLODwFpdx3+eDCAUdlqBDNGKkOP9Glm42B5ZtC
mp5VSRjBFSWA793IOAacxnyHkQw8mtBmKImWUb/iscNgZDffiNTLgqLoccF27KS5
97uqo3i66T+kq2HOUNynshZ2QGhCi1kyADGau7uyWzk1Pfr3zIkgP002u94rGcqQ
Hs1bWM1iBRWbPhhw8515uU+xT0sOXGDwVRSAkMxyHrDsQAtVzi4KlC00OJZ668/8
dYVXb7BSn/1cb3CLTtqaX9ymMQ9ftyr66SslHVNvRmBmMDrs85891+PdatMFk38p
Dcc28nWi8VuyxP0ULZ3rvMNlaBVT7afFd8jSWzMOBMzt/5BpS5vbbL1oBqYbYf19
bDXZZninVC9g1dGUO/EJ5BGZDpbLpt8xw9YGI5Z+Qo4slve7bF4WH+SXdtUDbleV
hhJlRzKfe3Dhzw2FfQiRi9XRU9eUehtVJ6ptG26lpA4pP8716VUYhmEOaw2UJNxv
1CF+RcxiteCkSjXJrlc5Sw/0uyBxceQVs1XCPdItQxhHFq2YDDyQO2e12kStg6qB
3UoK3lKhev5aSXCE18v5ZNsmzAEQ8gD++6sokdDKm7bj8ZX6cCArs/hINIb5db2a
FgzTKYLIS3WCwKKMPL1oEeae5i6BCu9vXmAbeQD5Mj8K/ZxztQ1QjuD60yMQmqhW
Lawnl3Ixfnl8OnfeQhNq9yXRjUrSS6o5z95XKwBo4qfdRCqoHbpoekBAZNY3GcHH
ASlRnOeJqOfmWmNcDDibCi6KuljtzkdjyzPdiXiOjss9lBQTiT4GR4SMjg+95X21
BXSRruTvAHTYV9ZtsbsNpFgdLvGVgc9HEeDbOnbsGX9bd8m6t6efyUGuI6Jxotsy
KA4+EAU+MwcsAwPvIyEiA1WogfExqynCLEbGclVgvZC6ZNLiOSAsW4PAwBO7qNsR
LuKb/ugdCLi4Ilf4S9yCQiUkYSaOXXFRnBYWvwOf6NhJohfP7qcuQBYp3ZlH4o6G
Zis/xzoE2QzP3MqworwwekjtutEvxuRne/0FajlJ/FurEdYJn7+UTOb55yUjRJyx
ygv6WLwizz8cniqxll7XEpdTxpu1OSL02YZvBLcRrY+25+T/73PxYr3AEU23zN/T
xuMjNg17vO3ZxBXLzrpiAv34qJJ100QkwQq1TOmEhnkPbYQj83NDhEBnsPIUiaas
AzXWknVWgVCCru5qeKNSbxr0nmUgXCJSQjSgMQ/FBKTqn0GejOqlc6Tl/v6hYiyh
kt8/i96dz9Mo3uKEGlws77Jg0iw8vLUA5PNU9whuPrFNyWjL5DI8DS8k7dqSLZD0
m4ROaA9lSYFVPeynCudXnbdWpMZM8ZAix+ZV6SOe3YBt/KXriRNxG28rLBs00ctU
o1VLuRdv7+gyK0O0gdwOx0ThPHe7ZyrKt4qPw7w3KqwcdiRF4VkO+KjVyC2JpQSp
tblnnBzhkT+zXYa1QmnUFRHbtxTQi0S2sG4DznQbIKs+r0UqEJ9HMRUzLUnOIlS/
BhEwcGzCSQVg6o1upk9E3+eu6ovKrFu0HyVYCP0+NTrIWBhRXlQCZwDjxlV/aYdv
DE5C5n0SE2GNkbqoRRQZ1g/sY981wseu+HqET1lnEI9IZ1qgXNYLw+etevuFKyyt
`protect END_PROTECTED
