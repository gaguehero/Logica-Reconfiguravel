`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9XOroGuq+3hJwZa/zJXGVgsrvdfFdjWfoz86Iog6oEfaNOt/Lk/LQCmOfSS0Bqjk
DRX72C0Ju0OvQc1g9BoGoJU8LTEVWFdaU4rhBf4I20gnIrCesdWaHe89C9xkuoQG
FKTmUYQBvePa1s1zc/09U8ZeHxKPzoOEJiXEeQTRqYtmfEp5Vrsp7eP8fK7U9VC6
XDJs2eht3whge4TeMvaSicUdU0rkijSgAyLCSCPEg9cIx1RBZ048UXdc9DUOPu8a
DYkFkJViPVIA6rTAxrBzHo/k4GFMD7ptYDeHKjIWRr/T3a4dFlXmWHjQwjJM4JC+
mCaN0Yp/bmOlo8+ZzApyAS25hWRnj87ywD4gL76vx0TWzWbdv6EQJF5w7k2Lf5rV
rgCHr1DF0SNqUTx6bgDGtkjbRBDxJ/fBY8CtFmFwwFFwrDBAQoBTWrNuPAarYiM4
Mq1pYVpHr1MK2QK5fGjEAK9JTVej1KTcTiEZHRItMY64On9MKoJhFc4Uyx/NaDWn
kYyA3sM/nLQXTmjRFjqIdmAS9Dd2M1ln7UMP22yeB9i0jBvmZwToJUiAUTaM8TC4
LyMd0WgiDO0HjOPtkPNts/HhWoz6MZiNapTOdnBnAfAQDT3wHjiJrg4JCdRpaMhN
O6liSYIKRXVlYeAfYa9fJYVtGw8rGk7ZjvjF9yRhHponk2X5fQx3qtP/ICYxhl8H
SrS+FnYqACa6i9frdRROJ4LA11ZMQLgfc28oWvkUGvU=
`protect END_PROTECTED
