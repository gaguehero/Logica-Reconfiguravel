`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WwAynr0CjgNvsIFnFk2Z2Tx8u9jaz5Lk1/PtjXMqCgssPn7wru5GRUNVcgQ+9R0m
HWW8LeCtZUyRjfM8alrL8FSYAEvwPdwgG0OmSG7OXncPtmBBMNcGv+oP53WIZC7o
TJQoNjPC6gBJDK3uA5UDK5jlp9dGV35qDKdoStFxYhb9+EI381V3t/+vd8bbXXZI
msYYWD/k+/bOD6fPrt54iV6lDPYSxgVy2EB5xGGQdtvuKTQ3A5dGKIJcdQiCZ1XI
VNa16Jla49lvKt8q7DcMWCZRZwMuHiJ4zT7eoTcNnRjE6pIPxR9a+xYGn5f16jUB
d0B6mlkq1E3Wnh7wjnQneDzdCmBt0MHx57pnr/cUe+JSteoQytpeR2c2P1laOQXb
dNhSrdgdH5cA/eeH3l/oaKh/vTKrfn1CJmhRSMWiuFLofMrZLVW4WEVkbF2N4q7t
jF2yAHWRrYa8GWMA7JQdS7rAL/q1FLRKy9ygXFJogwNY4LfefI2n3VjLK4aVNtka
GP6fKDbYkouWyjkO8TT/V04y+aIky6MFxh7KJPyrts57dlNbOz0a7utqpXx2KjWB
VPUkieThX9EhTIXis71m61WTcp8AmBlWUDPEKVqffy+9V9iip4hYJ4MXB5HHAfcx
WjXKtb+0lGFWt0ypv7hKEMAhqdy52A1E1ZxGevubYDFXHDY2VRPn1da51+RxJh5v
zJqASg48v0NDksFAKHlVRRM0crq/b9rw89IrPFrqCA9bY5nNuNpkDtJ84T2+0T3D
X8OllExDtJX6K/WmnEEGrnlsl4u9Zc7/ZiwwyxyBy69S52bgn+/wDCNUhlJ1TsHm
FAJ3KVNFg43dcu/MnMMSjuEEVIYtNwRTZfUVnNxo0CvRsjYHhUyI7tz9dgjWjPlI
in7bNS6O/r8NKcKsVmTUyBFxTm35hmlJD6e59kgTWNfkj5WiBLnYzA/1PQqhfJkK
gYmplgiUUDPqZbrpH4WJgZ463xikTX5bNuKjMY9erzhjaFpZDO6/Z/p+W18W9cDd
2RBs+p2SesNeGNsYidGNDG+4i+Nx0pFcP2cHS90yy8TrYlxUhxndSUMonpk/De3E
NAHiAxOpARdvTQgiH8sCYU8LER2klQ9Msk6nWABdw69Q3uZITg6wG8MaioTQGlgP
HgNCtse7A16+4N0wDMe5kmbFd6QXxG0K2Q0nTHPZZP9Wc16iwp4x5fT+VceEyjat
Jov3oBllmPWXNX6I9s47Lzsb58XTOIianaLi0UEKFGnxKwl2m7meJY3zlaiemzwc
Gl3oA4YMTefUBRfT3T9IxEFKNPtTZf9R76iaJCrvhvnZZxo5Mc28ApG75MW7h2Yg
tHZWnUZrDudRe27iyg9+N1YfU/MIXsR2Cj9AUtV9aI+AXh5LaJd+BpSG92xnPdcc
vwx4bq3oVz4hX2Q2D720zGB7WJzUIamNyR2lqDE++DF54ODPpPIw1YXln8GK8Mjb
8lLoBNHpPpquG/3anQ82/OySKV7Js5XkNE7ClQseivFDcBDaAFf1fRsD4LUW0Vfs
RF8LZN3gJ7gv+WRTTjEet1L3xqtaMdlhQJ3Tk1wKQKLjB9m3DjPiMmURbCYvQFpQ
NdPZl2uXEefgTki2ufjHAV9gqKcGxIUT+hHwixrnWcFwzlxkJhatVnPauj8nrioq
AEzFuS8NiX9802pNV//jK4CTsuHrYPW3E8U2VJGrDb5KxkKaLSi7zq3VomhNBTrO
v8hZWqDPnrLxSo0b9gUxNe6kKQIhXBSTsH352OHPA4mq4Ac8zJQTMGPOVY/IDfdR
g4Vvg1gvPnUiT82jK3y6n5qw08FhjPHlYkZkB12Gl8Y4IA48hsJiD2zUDYtJ5WPf
jq6tvR6nCD9xVCSs8K7r0RPqIDaSFsbnaId2WCvGf6r+hsyXeIKJvvsF+V/dobll
WMiqQJ6tW1VoorIf6dEPjreucOZZpKcYDCwm28ntVPQ7i1qQgrmQEJJo6/EVvw4D
oYcYy2BEfPxAy22KhyO2pg==
`protect END_PROTECTED
