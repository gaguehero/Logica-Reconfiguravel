`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JcObdiSxZ0Mcr0LgoOL71ODjnhHjMK8bANBTSztnuXGUC3QX699pG/bQmAfaNMuU
yfX4DM9+uWBp32TYX+PHBXfqkKoTCl+YKe5/RG87bjZPxX0PE8e5BYR1PDfeQN55
qi3F6redlr3L41t9cmrKuxiG+5GGdiCoU6W19Kq6Lr42j2ZAGmMSxgOy9EHGbCCH
kwvsxOrBqZGmj5UuN1HjIW38r8CELevDUf1x+3pn2XrKwxKwQS0UAx/HEeGxcMbl
ScTbwaTFdvGFzIijpefgClxwgyw9G9aWrNPP5nNGKS3iD0SNuSdTn2jMhosupNkj
a+3hGarpNpy6o9g64f2JrF2jjIbaD4dkw+vK+ROBsH49W6I5ypIxDuVR5F/QBQoF
cUfZ4qEK2bvgn7Q7ebSVwXnxRhNo54YJgik0HXP2x29FdsrbGQM7nOYwT5dXDdMV
h7e5n1ZBhy0/t5EjTf47XgK8oUr/UFp0WC6gWcwoNZ2i3IpqSLoUDrspwplH4Ymk
u/Zgj4MSftnihg5ER3vrLc6l157ClmspDj4t7ycORxil+5a7ayBoSwANl349rnK/
RxGNdnOXGpTilUwjvyFZKXzRnRYjNtn9S8BJYjWN99A4NuhQqrwss5lhGZIPhYFi
16bGYhDW/o48AqkEf9Z7JnCoZ7lYcJzlWHGdi18+zXauOBZ+qXaBCUxIb5QtZ6a6
mh6NAdqY9km/OyyH0g9k0AKKI9kmLm8kUTE/GoKiHa/8KFMdPnjpy6PbInzMCWX3
R71FYtqTxL1SEo5Hm92h3/iB7KZKTsxOFhrrUQiShUCIwnLz8kuw4e47T4IHPHHA
RYkWyoOI5O6yHIJ4ATA9HoT2ckY+UqmSyVGv0sMpwcUbNC/nlu66cVRKJ4jQHFke
cdW5rr47wwj2ogeXG2GW4sGJ/QIlOBTRtBRwhgT/UHmxhY3nyzigcLspmTEgxWC8
0pp5eclyTjj7626R0X7OgbHDQn56WWmwOwu+OjmY++1g5s2RG3L5pCeZUzoblHiQ
k9HEkuiUgGwi9ck5PyKcE6N0AdaxjHKYG3XRiVRPbcfGsQErV9kN9IXbwCwp0f5b
rlUcA+S3DKA3IhG+RE/N7l+X9bNEEo3sEwYrOz3+qk7o1/9+2ZxnwfqHm8J6yLZO
m+d3l2JB/iOX8n6dpgMvkkVDtG1DJ1Nvkno/TGpyxojja3ZJkQaBsG2zE5i6BoIm
FHtxPMrAgEAxX6A8udrga4CxIHVDJnkSkE+scpipqLI=
`protect END_PROTECTED
