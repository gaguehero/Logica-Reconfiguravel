// HostSystem_tb.v

// Generated using ACDS version 13.0sp1 232 at 2020.09.18.10:48:07

`timescale 1 ps / 1 ps
module HostSystem_tb (
	);

	wire    hostsystem_inst_clk_bfm_clk_clk;       // HostSystem_inst_clk_bfm:clk -> [HostSystem_inst:clk_clk, HostSystem_inst_reset_bfm:clk]
	wire    hostsystem_inst_reset_bfm_reset_reset; // HostSystem_inst_reset_bfm:reset -> HostSystem_inst:reset_reset_n

	HostSystem hostsystem_inst (
		.clk_clk       (hostsystem_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (hostsystem_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (25000000),
		.CLOCK_UNIT (1)
	) hostsystem_inst_clk_bfm (
		.clk (hostsystem_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) hostsystem_inst_reset_bfm (
		.reset (hostsystem_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (hostsystem_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
