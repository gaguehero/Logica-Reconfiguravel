`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/PIZW1/d618A1nBatoyiLW0iN3L6WxukMH/bEnmCHl4MxR/ExzFHwmcV/wxgkWn
Tie++vXyFXvF8Xy//lB/uByBNt5HZf5o8d3TkVsb90DWYCwEWQKXnyuukSJIfraM
YMqp7nkZ3oRNFVNRI7Zs3irGPIHRwSgrU+isjB9TW/9Y35+nHX2yzAaBTyNcf0j9
EgTQaggDcpu3COQ1nfekM4uxLkrkMPs+/WitoN9FfRRg4sB4O+pBwpZcaUIWe7C3
jFK29dWmpQgJ1Qh1jVXPcG5tdX29wQKhul+XT1S5ZIJ5Q6QRNtslOo+T2P8uGDWB
KkToc1mPsc8Y27VvMD6EhT5iNlKq7xQF0J7hk3owH/0IlZ6kZzzT3WYD+5SOk2ey
f48Rc56QCIPLK7NamWaeqZSF29VOg5jARq1m1sMjXVz76Ghr7Pf4iREsNJXfhpKe
ftqHQV8pVsMCvMdl520UUY7qYZ5vbbLiOU7z8QzwMO4zWlBofyj+fkor/lj4dWtx
A30rjAHBTBnirlz/UWGuwJy4P7sqrI+LlnpbizOAeBCC+flPwf8Ogzx1OciAJs2P
yyAN2M5qW9iyT00KXrrNo4HmNr5A4aYQL+5oKqwGJFra97tBhTKzd71a9Pv9Q6of
2GNkHvTml5GxRN+9hqZIeBkFpVKfDBgOsoDvza0rAXpqwkJ88TlXqVQBDSSd1nyw
PQcssPOjH3PGEon92JFL+hiaz0ZqLYkRE2Yy8vqjAEPQAzXJ/qTq1o1Ul86KS5SL
8Gnd6zqT8QPGduA+U/JQdCcFeuYmI+wZI84FiLaTb5pIMtOo7nHey3MlIsrDNCv3
RRPsVoT+AYIq7BOy8BeOJz/tVjjRfbDeUT80LjKcbYSnc6YT9G+3XDg/iIA4ux6y
OWvj78QndTwOYPR1J4SuscLcSGGzWFk5tqGAX4omRxN7FpeMZmWR7mL9Mn1uJvk1
MHp3NhGxrEEUBDFTLVESaRRZR81Uhz/cLz9Tem3Fk5cVe9RHVW830o29hL/e95zE
m7YzPH/8HXnvqjDPP0Bdxtmlkhr2CqJhaFiQ6PFuhtbbRu08rJXtkVnc0VsM4F5m
33KEV/tfilHNmMJrnGtaqB/r79nSylwWVuB1GIMcB2C9YsDo8LDJKiWQhHfBu1ki
viH2tqwTZicFyPk3mDCSsT+U3tA6da/YJ9EjwUpJw1GwH0Vxk01zDJEoQuvxG8a1
7JH5XvhN0rMeo50qk22THyPUm1qVVOWQ2urjjkOzKVpZOlXIKrE5BD85hTEhzTP3
izsV+0cXM0ARBW4GAeA3v92rQM/4pM3qjxf6bboqB+uQFH1uGb6sL0u0OX0Inkfm
1lTw/+IhkLnCM58Jul2eqUDdoHpTlDEXqToXak8GiHYad+gqQwi6UFUrhP99WxwP
a21xOb+ors4M4mn67D1PgQeIbtkwOAMnIH51VfiMCQv+xSK8BSpiEduLJrgvH/0Y
9ObkevNjNrBMkduR1bmHTieMrgILbWDSUydsqRbRlF5Pe4f+3T4N0yhD3PtR/QOv
doOzROss7TVfR2mkLSR4uRIEbiDWpXrl57pCgF1S26dl/Geec/ttY3biDJjT/x8g
RhJ6pp9RjvanWWziSVEAiAGj3Q7/oY+Bvm+1naHHcWq4iXfxNtP8mGQbeLFQcjn1
1BWJm/OjVRhOXWvPudK6zqDy8cSAPzVIeFFtcew4jv/c9BgnvhzwlghkpY8tyUv3
bf5X1beH9UhaDl2U76du2ko9VxSboW9zGH/sm1sO62J+qH6M4ZOiImTaT/jubfN+
QSBxa3ytenyyj+cqkjqQdVd6WlW4PKNkOdt+9bkxKCeU3iX9ZmXbFOHjkjA1hk3f
ndx/zqNDjlmT7Xbuh6Pq8oMk8xrkm9wYzxUNAIQHXSUeJKW1uBsoZ17dLknbiZhZ
Fg/X8S/zbJ1bCsagYjVSSlSq5D4G6jEBP6E7rzbq8rRmfh+dHblrtAVTOCavHWxv
iLnRRtp9Trvry/+CDR+cLackGwqchocQUPijUEAVPp070KanGDl1MQWFadl9V4Nk
PDhWB+/1dd+1Jb//0r7BZQ+RCYPsx1ZPtEWPDrV6dJwPiNmcRKCMg1fqrValjpCa
DyD63Jh+CqzIS0e6lN7vky2LizAayTWDaDsjHv7bBdM1yesfdmDQRttMIcI/KR1g
PjDm3F9Uj8LXDiwPAYCWpu3xTgB+xzza7iU4lPeMkGw5TZliW4nweBs3jVZm6Pvb
zIrcnyMbBCRY5mvB/fJKzIscMfS/N5anV408dtSfidzfTCTraNVmPZkrogrEZ0Qc
Qt5u3ZMCaNCuz94Qr0WniTMP5RbLR4XXxjAB5HEJvJwPsrulCCZR77XVCyC/KjJk
fJy9NncY6O7RyiE5TwS+xgrAzyG4jgc0Dg7ACAY5fF+qjNYEGizWP5CT2+za1gAW
IdseVLNHjrP42HyM7OP6DZijCPja6YNzon5d2aaKRv/leh34G1NAcO0FtoBru+B7
seICYqAz3aSilJpv6WpE9N6+Bp/yVfOukGaQi5+5VnJWutmL2wUEcE3DIUegEdvo
96khorOT83cYPdOVHr0Z4hWaaJjdQfj6OqDEyhH5iUBKygC4KN78cwGDoMuMC8pN
KHv8Y+7q2g3l7C/lTmcv+AJa/Vv5KFR2Ad8PcWEyEiTnl0/1rx6A9PunY0TSDJRw
kC2Ag1J8YIVnocv/KPdXdExS4Bqv610PC+rjxsyqKDwzJnBoDRMXpcAVcHHSt9W8
LgoRQDgLBg71YEZTCH5YseBSZ68DvA8/eJm1EVQXmvQzOoe02A1RxLSgu+5/gcXD
4zcV/PiBHB5z3yck7uWUQMc85miff8LS8rcCar9HaIBbM7ONp82aw2G+vyS097mT
EDB+9QYEfzgmcPi38dcHsYG8B43BbAshXAmNhK7RWAd/3ODoE4kykr6Ht+kxoEgs
hRbk55Yvm4VOzg1UtwaaXvsyVyMAjdrii4T2En2kimQYFaGoDNZcJUHKjb3aBJFL
1Did+Q7milaji/3xFuPxS65SOsSIgvjz6L64Y0czqWYsHKPNND0YQnddtFxBpKZO
SmBm8LVjiKpzjXDjs0YmxJiYC5sA+ZW1Yv7QknBLkr5Uc9HquyRWkr4pPv1urIKu
7TwB9N+eTwhQzUlqJHLtr2UR+djT/I0JqmVp3M5wV3Rzvh3dD5RER2roPv5ua9DS
Sajhefj7Y7c8xCUGQX1Le5EQB8n8CJKFetAd9Chul3KcnYKbASw5Zx2wt0YBgnH9
FNz5q6mT8NG52wit9P8wmWb0b+LBJ1BGKTeFV6gvfHzw/oS2wi+DX1swJy4hMMg0
j1vBYIq7bFhk9eIV4/8JeucgXv/9Dt3kymUSyTf7AIL9Kk2rcpmN/pN51hB/DwyP
f2M3fhzxx6RUrD/hbtT9Aodyhs/LKcdjaHxhZpxQHLwj5U/9FdD40DqDDPixPycw
aTqwM5wsGThtaIR9NVFB4leWWVUN99Sccy6LsW0euE4h9iZEDgB5ALx1deTomvYY
cMzeJIuqXBOHRt9lAVGZTLora2Il/Z7lnrOcORcRoISBijgh1ywHWNfkHVDOdUBb
gtK1y6S8sz1gugWrahAyfRtly/xNBJQ2iTGPWEsQfJel47Mowjpo9zjWe9xgGVe4
txnx7fGaOmgXA/9FQDtelgcxgJRWV/u7ieW8kvyAybcFNE97Vi56mYlvXjQ99jDu
ZC1iGppBteWllTNIsCfYk9lMIpxVPllaIFmmI7kBTDwJxOht+JOLuns4q4CtYYHB
ucSG8qF5BEm7rjSf6pAsfP1OequXUF5JyHgePBCOh3YHQqkj0ijnR2cUm9DLDYem
dWxCW0/34HJ+rv4P/alfh1QgzhRSNC7ZJXT/y0Tl63au4e2ohjJgBFFFOlTUk1EZ
+vKUqbMdYo1sM65TpOxXqYPeeEbaKWIS8NOoz3QR7n9dJ1exbfpYtmRUEO9RI4c1
kE5F99oHG0q5sauduFWNR/XBCDkKvHWmpKKarZy3GNy1YPZVjqBCPZJdIl0hPzHa
D8LGxOpJUSG/IpH2I5G00Wr7broi+QNHhJvXl1EH8xN3QvLQ5ULU9aq2M9CvB0ax
yuSEjA3n2sxLQz5hfI2CDoiMkSGbliJ+orzjsa0/vZ7lcK67Tz8dk7FxHAGnrxUY
4ZNYsip9iL3vjHEA1LI2vajXS1uksb0iWiaBDz1wU2NvCPsr19K2XlTKtDL/y81D
PZDtNAT8Qzhk9mAHGGLWLIkJUB6FlPvsXr8kZmHX2eJSIw6QQmMiRlHhm7lnYv8u
hqB1MALGsxlzNq4RiZA4lUCYaejkLS5OAnBy4pA0sEQyV1ewtIWChVAeaKrBUays
WeVzotwx+ziMOsHy6JPSIV1GRDqWNmANrShiV3r9NRPjzvMhovddL8wbMLSvgFuh
jtmyEXWSgIX2bD6EcGJwNMYG4Vju2nMGbtiv8Kuc+ArsGRMN/b6umUMmgrHIAp2r
1qSXJFQv872gwlEu+ZY8WngsdPUfw9mpcV9qlwyYFAr5ZjiRc3DXH2XrSCnIZ3wu
aO7yT36N7f5NGz9u7irsBuHCackIMEXV+r0aTfOuoavuCU08rrMOh1T9wX9pPdeW
s11r20eGwndyiX40EhZU7bjJJxIYgjEmQIdgEDRnF5lvVwWStbsJBq7BKBk8l3Rs
ZBNhrQlnv0usUm8QsZ6PRTbZyR4MvJ2gYizIy8NMvDGAndaUl6kZ/IUVKg+/4T6m
Hwco6L5agtuzIqUMEm21/x2tAxv6v2wYO7KUat8e1M/JR7eySbrKzoZKgOzQzTD3
P+xft+8l7THSxl+JlV9BOmT1jhZFgdtzTrqlt2nZ9cmaxg64DkOQwp64+zIotWW8
shOu1u5FKwCRz0w2PzNnys+VgJPdHHqL7mzf4bOUv4J3tpOOMZyxVfkWo4Rrrj3Q
h2dF/jSe9jGzHKDBzCvsygi9Hlivp+iA6b13muZQDAI33SJRpcpX2mC1lz/TjHV+
lGd+/RSelkm9p2LJ6Ecmw4WLbjsilXxnBUe3j4DZ1i23Tdx63KECM0pVnMR0C8/X
/dQVviPiH3oCWd7k+J8tZJZp7ZJwrYJE05jw601WUV35OV+CmYfeJsV9A1WiDX7D
jFNjb/GyXTCxUrwv4/5GLEoZR3quwg+ZwxoxECFgVsn6/U7PIJTK/na8bQZMYcKR
fiUl+uRCAqULVp6kUL0YR2QrCvlIly8ocvwrtuzwB+ODz/48mKtIAABNwi8DgGdq
AKj8LzmIhETcTwqbAaXqUHcwEaeRJa+HfpiuR+xKoXF1P53gML5EwMcd8yaNl8W4
0mFJPqhvUZG7AmHRpgWk0EcFPjigwuX7mon3eeJbc+69IWPvPsFkfYrPhBgFpjZ8
afNka/74K2GGABzY+tIXCaG6OJTXWQGa3VWnj3OkfPHx670544wGUANLEH2vGL8C
RMC45ii+VKdldP/MGF2ObvaHlt1xK7+RyPRQbL/jBz3sYge4VBthfsZIXyoc4D4i
uQ1w9H6FHvjt3NJpbBgJAR2/lvNF5XxFbTdtXckTfwUI1PwggBJw2cERTudJSOib
ei3IgzNtuZ+xuroBZ9f4PiR3z/XJGqZiwOb8bcnB+X+jyGOofhgWDfcEi96LQKmt
+vhwX19ZtKMcGGDNztcccdZh4n6+lq27OQu131MfiDvc9+162dr68rkLzX0Jrnaz
U//VM6mbyg5O8+OON5D9Q2S9hLxR70ZcWGVZ/hlDZZofIpzMChYJNMfA8Ocs2aC8
eqOZ+McsHrkSeZZZfNBajB9ziuLIr/zO8XxPF9BNhK5ccPuA0IYFBdTm0ZiONDSf
n2MBGDWuSJQyjNOJCsnuqmduwzlGCkX5ZLyv+fhY82kUx/rRcAuS1aGHZX4Tp9Uu
xbh4flEzq8uzy1Np+Yz4YPwgChPS3m/IJWt/AneSeWjsyLCbwSkzgt4QZYsOSvRm
OqC9sj/kfKe9Xso5EGpsqyL2TW2JYNC2B1GU84yXfdOX9jyWdZl7O97CV32T55Ez
jkuQYa2T+q28MP1LXG9E8A/4rhxCzDGDW73Br6N7nAzuf+4qPKVbBfFUGYmSteHc
SVVwzHapUGArZrZBKw+MOjbsErEki76C4ZYnh5IgNSbQvo9J8/4rxAasjTqvcqGY
J/naTeFuySv4Nfq6yA0s28J7b3HJJIh1FMBz1xfYU6iJwGut4/JfhuCWc2m6LCgK
lF5dsZg7TIIqJD1pFHqoH3dbOwPGjhf5IzHw+dJHgj9IOw9fO3PB/0+LGUxaYkPt
EZDKkule5pgHgu/AdvQqLHRcbviz+jjgG9s/A3FDMETuquSptEiLytYU00l+8hYU
0RPjqOVENCWWf6CMhwbZx4zpa4H7QF/lt+lk19k9ZwTCFeX/Y8V8QxprYToPvlrm
0S6W2eLcU+X0PpoEK3rZ1pLBa+lbDhiMci6U36nNUrspoodMTvvpOdM/3n/p+4R3
nQY7roavGh4gsDxt0i+AhKbI8bXNUpeYLmBVncDijCVViXxVaNqc5VXPRjM+d6Cs
BxvthMNHtcN0ovE2np/4vfhld/H0ztRkhQlti8WJp2lUSR61ZSqQnVcU2re1YNpU
w/x8xbWYZ0tbK6kqKnkszIRRzrEc+E98sUfldRaRHyrs7q3x8RRxuKE402TXyah8
HSUsYP2uL6fjH2SI69TLRaqmVluUP1CF7uqw4ERBP19YLF5jWmoQnOEp5fJ9tt7J
PtFsTZUVy3jo0hEUNAKBXotpLl1h3t+l+raS8KJLXbGOcxsvEnh9RRfOfxvvBxQU
c18UotC3+kfv9ApgrMLcDVFyswurs4HabS6FFUQwspMyiel2EAICe93ZY8RLRsQT
niy9VvJixJq708t7WmMEqGFQYDzhOW1pHxCWaSYLeEzaVaywOGNpdyiCOBBHtp9r
pl2ZdfRYBp/CL4U972fytVZIucqHR3jIW11Ivj/gZ32yxGnqSwgr8xgF84xdNKtN
5XOW1w0YT7kc1vlxxIBlFKRHVmpvBz1WWwox/UxSf3XjhvBFoWsNKI6jHb/K05B+
QNQ1aERMU/UGUwlc+MJjaOEX3gs+GGD1DQq9zPz8nHhNn/bcn6r/NuK4otlHG7R2
Im1aukyEotw/KojO4JVDvDBwzHP0SlT53f31R+JB3gInIbLFOwqa/WoUq90MVgmt
VAuSKLmA7V1BLvSeONL2zbyUzCalPNPnAcrkkX+w9U/nC0WcdQm54IsiJ9dRTrtm
LbCUDeMv6+91OFZmaCf6VjnulkoqWrSCr1I5Ffr9fOoJyccMNHWjA0apTrjsNy4r
YbQZjivHI8b9M4T8lrKqQY0dXoJLs8fHz+dgp2akOCryDtt/AZajpI6yjeiFjQ/B
KorLqR1Rb3yIox3oBxSd7oIE0COuYrY//SBZMivEL8IP+hcSFqlN+k+QmPpYcsk1
5W60pCD3jCWGcgvjRi5S9PJysdsJSlPTp1fBDHf4Ao6UQ0InMIsgp6cxUKLK0Rew
zKZ2CFfQ46gMY1nfbI0Mwy3qMN9bynqMDys4dgtEF8mEXQQtR5I26N0OrB1kwsG4
TnJjNRuXVlA3UJrBn6RkU/U5ulTZmiBlIBgomMRYF/dJ9XeMBCdDnVHYvbGZKSdL
Y8Gss1qhUnTXVrt21e02powwYJDYnuvLYYGFH0aOilXZDWf/arOxSfMKUoGlK85p
`protect END_PROTECTED
