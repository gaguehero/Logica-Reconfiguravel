`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwevRkRn9A9AvafDLOhebd8JIoeqYtV2fJeKZ8A2WetCQZE+C/Y+9uhkZ+dWYFJ5
FxYpimSa18iCeVYjjGeb8jY8l9eoEOTcWnk3YCKuHk3JYAGZcXtuu9SylmBgRY/E
LFLgNwZTLcV45tNQPe1aRDNf7gJg2zoBqTgj2xPJBcaQ6VNJln6IEjRlWXIRTX5j
OWgKXvQvcddSpGXYoolnvLqT503tVLCUDDX/PFv8xqQjiq588JXgf2CtU4vRethR
s8DAXbGMLKjjniW5rJLbV2yJ0q3sGOdJu4FuR63ebEFnKSbspuiLzWXi45h/LGLf
k/ixBIozgYnTSdUGvGpfhiqz/mmwIxYBOByEX4dBchwAQHxT6/+B5f73u2/SsypW
cZ96wSfHq1UIRt38HaLdPQqb3RjJpYR26+WuHwJ76HlNXS8w4Hi5Cjpqf6F4Xvzp
OCqya4bh11kIn3ehJ8ABi70+UB+xZ8zHHU6Jpxo0SJbAaRTOMYrls8G5OuN0XRTh
fjmsrdej7+mmcr3hcrV0Esa1anptPg9Hsj1yubDejwZtkiNqYOwEIfuBFZ+oW3ol
KeCdo5Md7+8GRqGJlSdLuMKYIUJdyx4xWh4xBX+So9GdvDFHUJuOK9V9V224hTLO
c7UL4DvvNh6PTLrKuqrxg55sVVYwZJqmluvw+38GiLgYZ3pAbRd0De3mgWQ2iuXX
Unm6IrDayfsePldB2JAV+y2o8fktiJ8EzRvA2LiEzZV1Q4BEtmdBAoLxGh3cCnmc
5ghb/L32slUEQ1JjawM5SzbMIL+ZuDjz4pDqTLgWNcJ1v/hkFGHT2qvkKE+oGP46
QVkrGNGYu3qAiy0dQkNtFB2HWiu7mmPWMBeslzzY8e36Z+WfVv0yHqAVj6pgoodq
5d2mc2SCc4CrighvbhiQOyS/25fyX+rdCisIqPaS2Zd0r3vaeeaCMc/bPlMGUpt5
lyx5Ya+BDwymHz+qQrNQF4pdDygn5WXgKlOnk39IhWtkVwlmSza2o8a8TXdrhKy+
cn+o/XRWrZ8HDLjK0J0xH266FhUEG1r0snNMay/DV5E3cvvLC6AeeEy0nPWsK3cI
saPEo6lUzwhixbwU40IZ4sQ9Qz34qEVu78itfafAFnrerkQmOyR5Sn+EL3/c6i/n
z0hiVOV7YiDcSsr5Q2uCUqTcFxb/4s17OHSagF0wY8nNhXtK2MdeYtY7sLAE27nU
+ukLmDuX51zgJe3cMsusSqpmbbh5k2kWH9J+Ui5wu90Q/pPF9lvXg4jC80dkrjgp
jQBOdV+3QlBf5PbE5c6UfGCq+NwMqIZBpqWxgEbT7ICUJXpWFovdWGLXCJvqHXeZ
zOXNRyiUoAViI92fQ10WPVWnwj76UhPdnufcWRw5BOdDeBMa0/hRGn6f37SkbaSW
U6Lau4HcNSbp6oA6sdu/bepF8W13IF7G8v0bnM1X/qApJK9X2VZjma6upa1cfYVW
nSxBYhSwj2HjYdrJ7TZX5KUREGA5vlCv5zt51Vm7WzMzC5OMPx3NVbCk+n6RgaQZ
Z2oK+wZc7SoUziiuAvuko5aoXoDcaGS/cw9qHm4L03rHRz40j87mhfsW5yoNXI0I
//TgBI5hQAQ6CQxpNkHqk76HqHiX1xCQZVErO8ONz28SlScQ82fuaQUzphDFO+5Y
Pib4eW32cbWmiOS1Odxy3CV5+eaxSlu8M/Dlgdw/o3etABsrr+BqeF5dCl0wW/eS
NGuUQoMyK0Ry3FtCW0vgZYRm6yGT3fhQro4CtiktgWU2QDaKCJGcqZyl11VA0Pwe
w3R9hfy0MtwcWCE0pzDMvtYDWLO9Bs8FDjpKrEz3IVSOGWAGrGO5XCZdhNSi+bdb
wcyzQEt9sotpoPthCdnPHpZE6kfZ7F1PFDsxgyGBuWE2ay0biZqTHgFR62MdKziE
1vxZ5J3ukB1KCK9F8GwkIWE04EmxzgQ+cDeJX6C9HIE60qztec5GmYFftR8mkMeJ
XWEcPfOJSAeyRD7ebobxFOVQ5gyFo0BwHLJBwJ4xQ5jmxf1DMPN+W/prO6xtfm0x
`protect END_PROTECTED
