`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BrA3nkKokjFBGb+hKmCGc3SQ6zX2JFyIRlaGlNlt1dq23jrKXZwZY1jRcd5Iuo6N
rbtG7m7mMZ2CDPnxRXVUJlebK05Ntu+1z5LoL3ckWoz4276G+M91w1FwGBDTVoat
HUrRm/r/POFgeI156Xd8HHWLEKZIOO9zaGh8h1BCqHx2jTHTfVoejCytZ0qQ93fP
e8ca6OMkHoOu7dV2W7V13YPF3oagGMJ6O2x1G6Pnjv/RRSFsXZmIBGvZYY0Utn8N
Ti5WUl5YbF4cSpmCrl/KmmZNOHNEUHNoEbI9+0yQpO3b0SlbAmX9huSOP2dpX9JY
ATo4oq7fHRbYNOwUtTIqQAmOgniOHx0JngOi0IMpGCtP6Ub8Bw/jH0aNLxuPusBQ
yIErixLIOSUYza0S3AMDoFs5WzZ+uZYCv5zLCuPMZYT4xXY41Sm8vVPwFLg0xjJz
b2FIvd8zUSd6yuE7gupTaP4Uir6kKsR2u1y1T9tXsnfkoa4+i5JxVi6rTEUDk6ew
drdhw8RPUmJf7E4MNVxf6EPBvilZ62M6sYhDughpKS+7GHIog+LST9Nf7AZGLrjb
yiG9IN5avBNvyOm6xxBRt5+VyzI4BAQ1QcygxACglYSc3yutbBJ292jGc3kc4M0z
0jorwk/Kiyx9PwzzixBjWe+3LRFYfs6u96EqekuC7jBkHC81a4cGZETBP4abdHyT
Sm0016ettRk3l5H54tr9s0++E3Tii4C2s1YWmYkb919NE4NvGiJhWFdMiqfPYA1U
n1tCnRXs0CUrZpbzdbLHGuXgxn3luziLXKr7QoI5n/97xPWI+EruJ7vRVEnLK3OJ
XKxQcG8J8M9DmVkkGd8nXKDoP2IB4bDvJ/6+htEJmXgyOc89xDhCPC7QBGSlFx3p
xpmFKsUAPWvc0RQ+cJ8IhNvyF1KgFZOyaQ6wIaWfxj5ratlxyKagQWVqW2SROTAC
SqhamRqEUKvCCBLa7WoPgB3IJCdX1NWzfj7IPKTC6NLc45ye09AUf2a03D4ec0yQ
vfiMtnHMe+XvFLbQtucz1Hea29PcTBZi21cs4g0Tx1Yp+MPf+NzNollaMR6zcYyx
A+qfAj8I3Sk9vzMBlHpvHZAi2DImP+6a8/dosKFmmYAnAXkLhA3c/9YFhO0LBPuD
EdmBXxwTJpvP/n6vRUrFhRICg8dZ+yLty0ItplOxQ0dJ30iWjAoGrBwcKxm6zH3n
3vP+oJ6YhXhxf7n+CYk0l4NmDYg07XFfZbopszSGg6y69uikzUMfEJpoiILbQCIG
ZBBKfDvvlHHUDenNp8ZTqm4Wb7Q8yzQeoJcRGAMMtvfDzwofjBrwLk8wuqFL7h6n
J3ROhFYfKCRpeS6dlbuoz8fXvrvYE1bW/qMgCXI0K5ThW4D0m1NW3UEryiDORVpk
6XFqoN7i+8VkMBxgq7/CohS6PnBT7s95ZEzqXjzY1wVGUEg+E+ygRnl8JBazY8sZ
vdc6WONxBnWIq8ysVGUvUnLPuqDpYeEgoYYw019sHDTl4wLA7aJHxnMSxqWN0J6w
iqif2J1wY+F6TuV0uMWekpjAUmpNj5enbiFKeURQf/gVJ6pV8wEExYfPGkMp17de
fAhlTML7MoaVhhSCWpPHZZc7DbM7V19ZDcXqfl37/Qwq4gHHdZRHc27tMnPIH/P8
9HfLnSMNHyes41wy/+RL1RdmvasRKsJnFA/hrLuKjnSQyNE/4YbX1giV7dOtdMIH
hjXkTIL8N1HqXBhd+8Vmpxpmi5qG3SYSsOWSQ0Yw2XNshPi8bmbXdDHj2+xEVUG7
rLzmNfkpwss4RUBOZ178sFPFIEfhEOOe17EWmyxxIZ1yOoR7hPP7IydjeivVBlLT
5su++a01CvnsCi5LupSoSEMFftKSEQFc6jkt8fZG2VYuyLAlFnBGZo0rcv3gNxxv
bZU1udaA7t7XFEU30nGeSbl+a5u94/zo6dchcpvI1t3gjrdAghEvw2YMYOE19VBg
oRSXiuVeZWKFLH5X4iNw3mpbWTs437KhXqK8WB4YisnVTeB/shFro3YEJhjVpljS
iwo3jp5zQGJL5EFcj6jEmKoE5Iw0XKwOMYXw7uMTZ/VLMKwlQcTRN4g1GR7aTiRo
969bbxMWq8+6AmEQ7LpwmXLtdTn62MGTywuMqbAMxs575XtV30FnmYfSNcI42QR/
5u5Z6H7/hOFqCLYv4S95LtuGKKp13A7soMGFpTiWQG6d4HoBm8RO7YxPhghcvYfa
ROJf4CfPJmN5RVbxYtZFztYqndO4GvfoHB9j7In/YZ1HxePaiON3/lbC9xPKOP4u
vw2asn6uSuI+dwCjRXgeGorVJkqAY3aLLZnCSkrnE3TW0UaswmyzyaAMr5xqli3d
yevQQUqlFnxrdVXmo5k0EEL4jmREqMT9tQYWTrsFXPAOrR0je1xbA2/oQmvNFmLH
MRfN1CjEWtNHRgHiOyChpp57SPosZC4pamumrORb0/TWPo7AJXGK1dWu1Q+aanR9
/b1RbUpX9Wn3SLKW4Nmy0RM4APOJ/DgpEWUYqwDYrKq/NoJzpqnvldgRPTOMLk+n
gwrsWeVwP93O4VAdQFmbJ+UC/jDxZ0kYkHWXiqU8xLm/yUbdzol7akELbxsMh6Vd
hPws8A76BARwS+XjHh3HE/NDgPsWy6VgK0WLQHvaMIRvJsSTcKa/LZLwhqLB8JkW
MrAevr+lAAd1lBU+SIThZI+LAVJ3dYtq0zpCRy7kSgFDOihh/Buo/O4SpHz/zCCD
DvQ24qLQzw6tydWSx9UXZi8O7ypG6aJpJrLF5kiNFjqt8x/akA93ZRcx5h28rDvn
3WhxePHhXFfJYz99AOgFgmH2yb68tftbGJq/RUCGpZFkYuUK7g3NiqtZeAwqMof6
IuOS3EGlnRfO/We7enQCklvGy24ACktisfsJNtfVJAHxFpDXNYF8miLJ8UMQqP48
PYI3inqteOSBMW/rchUFLbAdCmjYjYdBix9tKRR0hC8FdGsquhfi9npET9bPHKIf
Jdxha2242lQe/nBPSxRZ9y7bcdLIGs3dLkfeheCu1rXhDgq7BMZ3FwSghvt13Td4
DSYloJ8VVDmzihi0fLHSvsa0d+HN/oZ/LTeln/KzL3WZrpePRBXIlRWlJqpeuaB0
7JzLRRP909q+X7Md2HpUBJLnIE5OknqwkxbADcVQ38yv6rJKMVFHIeTNTA/kgN6N
++c0lXUrJ7M9Vuc1iBqUXP5PwhVKwwHtbLisOkRxX+Wp3g/+xyh87iAqLh7U8yBi
c8eUpLR0fF8Gn7gCISejn9tgN9+xLbrX+iM+uKhs0++L7j4Gw0+5pRRP00WbxjUL
M4aKT/3IWRZIY/Sbv+641DbpWULL7+75LzswhfU58YTaADGSyoYd6Aq9jsupOudc
TtUYfsZabBiwCVh4S3POSoA1QrEkkHJFBDMC8lbjwKIENw6v/0+qw04bAwiThYBv
l5xAsrIIhqmvjLPK8r54altaewsOLOsrPOQcUbGWk4sF9Xl4EJ6wbpC5Wpu2L8OZ
louqIsYcqPo745L2H5uQj2AL+7df1yWHqUtMXJwws2PHunmRH7/Itq3OTulljdKV
+aoB97Q64P9IzXWS5xrO6hh1wguZuMA0wEMHqZ6/Yyb9CtzKccYCe30pI3/06Nie
MEqtQoKonqYcsnkph43I8Chr2PpTnqdoaMi3Zo9ps/+4OTmZuzzwTBPOgsE6GkVv
8q38XINRsotsW/rTNfT3UMzSfOLNYeXeyctudLpqUX75EPqOslokIPTaZyn+nS19
TpQT0HI0UUlMFoscvVlM7wb/66EaZKNx76LYJk7Y53vBomnX8faFUjlfYOidngyN
GG60Yv2/5tkpGBLn+RaC5A77DAl1t5YEogLsNPESLKNLHOy6n/ZfbZcRAsVlInZp
BmXetrESvs1qX3Xy29KyL6hkDawJZ9TrQ/M/NeX8u3UladK640WVzZCqAG+OSfs5
oPBKBfwuu8+bTU69kNK0j/eQPBzW4Dc+y1OwWRTkCEpEmZpQMELRWfA4WejSjJb7
Y2opi7FO5idDrF14zVPAviKV6gVeEc/22VQjgtNvxVX/Wk6g+gSP5QAeYBoxn8aM
b0rLeiPmaWyGxt+fLCnmHt8Un9bigbDt1JXcvFIkMZjRMjLRUpXSdffzMAf6mBFN
Fdfa1Wfgn2GAlP3SSzeuH6pxr7SjVqn2M17WNIMPyIz4UZyAx0TwEJ71rkOCDxX+
HT/3ZLSio4HjBZ2Ux5Ely4omp1+qOJU1FbCX6N1DTpJSqafKqRaV2jbU8OOTc566
QGnQjofZfaT+c+IY5p9UlqmoEX1yBozGL1aL6k7fhK6TFt3QO/hPdge6kq3EWdBl
1H4QcW3PPBXvAKT07hwVf8fYnyohyUSGRY+X+kB0VCDU3oBhGnDcBsLzSn3BkW24
VdG6pLm2EbHhN4za5D+kMeGqAvL0uEZcSlc7pjbDSLEw76zoUm/O9IrNJQChWd3a
b0TmIlAoz0oObbBai/C8+CeeIyXqZlc3rg+Wxzj41dKfV7PE1nG2uUZo0aa7jBZP
58RMT9/XZfABxpwrszQGBdzSBR/O9/F+UEC4kMqhdseyWmYSUfdPaEnhnybyDJcF
ndGyp76rHWv4qFHWwvDhjTyUytpLrO7374p4lSdL5IFkDoGYQ5w9geT+JjjIOjfn
82jDXOwaWM4HPwsujc3QFQfYzlE9Nit1pimTYVEC8WSf1p1RgR05icA8NoKcXiRH
Skpt/K0tzgVppI3I5NoMpem0MOx5zzbywOovU7DQ5+f3M/a92bXnjFPKoKsXMY+k
mVmm9IDOvjSkWu0uqUV+anwlJW821hfm2jCrXKDzj/XGjLTHmRoQ/1QocnaiEOX5
PTOzk+nsL6fatq/XxF4ls5CqqyJYKOv10mRredOIOJLa4TpIqYu2pDSfmmUNUv0J
SqLJe77goa4g/1EkZ7pxgTGbwnDqCwh3QzpQDbFffuh1Zd1RC8a6Z6kEXySWi1NR
hD35dYhZXhTh7dsrpX3/Nqv54BM9bxwfK6OplRlBu7HuoS4mHDQPsB18v0QduaM1
ObyWDnIX2QPP0mnpGdSEO8IiJ7zcJD9eG2oancjp/z98gKskVQyw+U/T5+sH44Z6
0wvGO7XKV70zjpee2bSnleODq0kx3HJmWcN0UQtqC3svcl8N9Opr9ty3Jg74hku1
aa4QZytucFwxDwQdbl0c1Y9B3WNKQ5RguzfmDLuW6+J6xFO3Oom+InQi+pqwn5ik
+u4hTaOob55siZQ42pWxf9/KSTj/gFW9toKK9LKrHXQfoqkBwkHcBSYimCHS/tmB
uhUqEeFxqC3put58CLW2RAkhT7CBXTBFjHxLPj9M/fHpKJPkHvo+Ti6pwzjus3o/
9tgHlCCqCzVqOeeCwVRS5nOvuPv2yiJQ3+tJrfok6VogyJi/maE8dxfS7WJ8/r1C
xCDyxLedYFMXq6fCwaP2+tu0KdMeqDp97LMmR+tfCxOEBIMukAB/+pWcDaG9h0nW
VMZ6764M4Z4Kjblzs2JWbnCXzp0f9W/K/+Cl79R1/4mytE59eAdEzCzQQORkPN6c
8nhi9FBVlMAtAX1m2XU3JXMG85ig1wUgK23VYci+ERH3EotWQzJSueN7G2ugC+NB
x+ezZPawFb21TikYNTLWo1XHVL60f5IIENo7IsZthkN0gZsjImTdy9263oybVWYk
ZzlyQcZxc6JyVgH8WmnGBnnRmMaBjB92EiTkKmpLwbd6I5kwgXToggXqQt7dn4U8
n7oePMZuf393gsVoeYmtB8o1+0PiLGcgAkNq2xCw+FKTKIoBL9+Eduq+clBtdovd
wraRspDhTwKq6XfLUnWSeHVBxCJmL1LW0PsylY/VsWZnFNetWUn0d6LcLR1KzEw4
IzvmaSNdsT4IbhzU7aYGAM44UsndEMHcYfzH9wsY0nQ8Aatw0PdvCY0qU8KaeKxm
9SW3DLSRPON61g83qFzGmUuT4Di47V/JavWAduzsadhLTVqVaMmoqz3kWpfssYOc
OE0XiGCOon80uvbV9llO12BsedoVV9MelSPYRYszynpuGpqTw/8KYIn27feDOb0n
T9enUXmN39saYl6WQJx/3VlQznaEp03NpP62DDNd3ctCQQ0IRQqeze7DmRTGXU3i
Mu0lr0R3ktzuuhipoywA6vnU1B+sVV1rGlQRq5Vn+D8fV8e+SpLxKsgbSbGI0keE
zGwgYcC8SzetsVeQ0mPcaj78wi/0LCy/HNSbDmKZ36xnzmL9Ycj7VRt6cLv8AjkA
V0Q2Vz2k30oWvG1k0/eA1S+XqVVV6A6BHBPT+EkZnFiT22KAXYWfpY4YoXwmMyEr
XeGqY7SmqsAIYAQh/uVfzvpmNsdTWpTnvJk4qCSCRr/PALoi12qivUmqNH4Nrxlg
RRZuFr4Bf7w2Rmr1mo7FWgok/qt0I65dB4cjsn0lLFIRGrHcgxTn16GkoP/x+ogc
bUmg0zR+uMbr5o7hCd+Lc/wU/TLGVBx0Wtz/M+UjyMA2mIOs6xUiHjNVRijh+nzr
NFHGglE3z8ANUsoouQkuq1UOczODxkirIi2TWntKlMgrcM47d02E1bGpxpWsWB1F
gZNyEfUa8lX2LRC8VXuKOBr08Qq1FL/hqzqGVZwp6cRdPlVWOBa40zC4Sww9FVZH
Hv58Yun65TiLJzJJHwMftCVMNg4LRtAnve9byktGOez/pXsaOAqCmT4mXlERvFC7
IjLyo2QFrFO5LdTaV7EfiMdlTN4CQFvpZqceBuhehCZoPBUVB13XpTz3dpSsqHxx
HssWp57L0j3CEt/p6mC0vh53BWWQWuCC4RK8C1XwYPVkA16eVF97l3H+BYY64Re+
Noj/5Gbh3xoDABny7ivWeH76XfCwwChcONni4l8cekRWSTjJYNCnPGxA9d8Zr3tk
ag7geu87HRHvNbfYMYsa+SfroHlXjwbDDgo/iEuKQoqy46WmZpwiRXu6MnG+Ci3l
jlGcveLswOJ8vDy5EOe6FPZWIMl1djgue3S7/ML5ofJZof0FutTLeVd5uGzbsZNO
nl82T86ijRIxepCCcP+E0V0/oZRy4uHZVCbfa/dNN6ADCVP4MMMby5Z2Nn86rjWw
eUmnezMRCc9QvaOtHaDwa5aEqFoay9jCJLPm7RRWcisr7ay878Cs7WNelf6MQ8/T
ERzuTW54/2d6ebpiuUJ5cczjaJ0n/KduhouJNExo1ABCCHG1wlO4BRinvDXfmWCJ
NqB6dGuu42Lcy26FfyDJ1C2g+pKsGYp6d0oRuDmZzSw4Nwb8nKd9WM0eD5OD1n3G
+I3ic3UyA3A+ZcvVNVrMmOvafakkyMzrN28/6oAOj6hSz2gvaSXzeB0Tf2798TCt
ZUfWPI2MJthO4v68eQrjrZtEA4p2Qi9qsraPUPElv0rMj562ZlBRGMxu2J47z0+I
BVp8h5r1i7GJRnCAqgSlcHjkzyfJT7wYGcb5ZikLI/l2lR1l6lbqaLn9tvuKOGs+
W2wZjDxulXhjx+oP+Mu5YqVHnZQUbzWyccZyt/gPIZEvKuXCBPqxYNWLtOWw5UPS
JUsTCRDWwBeTL4TDzxOiYk9hmxdPSa5gKsSLnkF8HSEkF8rogvsb9Z0bA/CCbNU3
v7WPm4t+kqigMENqHkQ5ym2v2k7rynhM73LssQXEkn0Wqq22iINRi//7aTU9inCg
PEwrbyNMMaxIzWCTqZ1Uahpkxjm0HP3LGItqbTJOjiOmnebP8lLenNiexB9Tl4sT
Zt+j5daj5UZQzTWpbtoO2CPDLHI+6i55TSbMRifTjJiR4VGIzmnW7Y12WeSRAlom
whTMOIGXlFRci0jpJD+C5pqSuwiPByWnwU/USMntUYQ9P9AfwqvLbUZaqTLBNk7P
2Wmye2u9ZNpSYxGxUZVTXHeQEZ1RU8B1AApFGw4bj+cNTIlktMdJRA+FIPAuWsl/
pCdVi5ktTh7jL+LHfqJGI7Y3b+TslVA4WgY6+haeiAxaqlMIF/VWw9FKS6ABabql
73cTkhRX/rp0WG8EifrXD6DF5qm+5V/CC27/ki8sx7W3M4EJpFlMSsjURrOsqIu9
azPYvE8S1RnbufZoO4mcyHsdWPOBK35wGDlN3putYGWbgPk6FLbVFC56fBGRqK5k
J3t5EcnoqB3PkrqwK99CDad089IBJzRZe5LYNdR56aPvQM/2WkNCqAur7f7K7Fbc
ATT4K3mXLFgjDOL4TxwvlA/WUzj/snC9CtmFbaGRHPb8FpGNkNPPUXmsid/p4kMv
OThiTQzcDta2Pcb/hmMzVg/i586+z34pLMYngrMnQKVfUzqYH9IJ4qL1cjIqlAmt
TgT8Y5RBqbhg8wqMmBuuEWsWxN4iValqSDARIQ4JNF4N9H84dQiw8uDfng4f7Lpl
l+977GPfMHy5snrUPIZxC/L4dOYbNMC+zI5uAhHabVnY/osdKG0Ev8PwFu5AMku9
UCO+IHBuorJHLubWjn2sCJz2JqWZ0ELAc9GiaEFSixm0/FBB9NzOit14SDLxTmvg
3GxCMUDMRG7Cgn5ihpjAeu+YClXB8J5U/8euW/qfcUTPyIW8YtOe72BkLu8VkFuH
ZU+dBTVUAHpi/pPGYF4rgo2FYZXH974cYBptXRUbtZUYc+Gh+WfHyrUx/LBYpBDS
aIdEqQmqtBZYeV2xQYAg30r083D1GK422JoRY8LD9UR0+DNyzbtDvEpl+wuNZbxw
7g3RI17WtsBeQt62smHe4gkf29cACxTJUOxuVp/RfakqFv3XpbZROHigvPuXKZon
JRohbPdeT8TU3HoSd0AL1NYWjpNKMDfduPlCG40uEaNC60P4BWf0VxAG8XMI1mNe
n0S8YaPG+pN9mtY5Do/bQ3QxG3yYyi/3Kt/9YfplLp2oi3DUJVrzgBhLbn4H344G
kOILCeCm2zShQ/fnGC24i7gm9p1+Euf3AT3gjAsguyE=
`protect END_PROTECTED
