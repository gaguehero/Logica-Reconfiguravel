`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XemFigffmYeS2HkBU9iVcH8zHi4bEdFccAgRw+F1H5vTNwZyugWP5AvYblcvBpT7
1YSyzo+dJaSDALGoT7LBFOFZA1MdPLUlQscBuaXecJVmHPpA+hOIY+hEpCAs8kQw
Wu1unAqlTN2L/56vzhsoG1b/uLtKYTROzhICG0pP733rKlJzAedp8FwIcRb6Bglp
5PQfGnWc5U22nUaFtaO2eoTS9S7R/rtnmwzGQwQ3tuU5j21U1L7PBb/EGsJ/jhqB
Y1J8v4YvzSGKbB6fPPJ8sSLbsoP5KyBBTgKXs6xtkW/mg1ZNSdpv+TydqGZ/+6hj
lEdcTF6grgAFv/DHapcT/hFZIFlj6CXVTOnnxyek0QCRhFUDC2xuDKAO7OL/kdf7
mGKGwonZR+TS15VxZt8Fwe8WSIdG+oY6cRNjrpj0gL/n68s74QTnAFUJE7xpNE9K
3veDtUye/+CsACAlc3bGvT+OSahKtvz92Es/SEFoIlFp2yagcaZ9eQn6+CizpCUl
ArGn9cygHanWfGoExI+fM2N9mGn3Q0CaE+L5Psrdj203pLWMy75R+1mlSi2w55PB
tt8Sga55Ny2yrPYeLAaOwjN6mGvGsEk7W9jai0aE9FBs5ekzquCikevPWkYSfuK1
L+G/GsqzWJ20fqETj+01n87Ja6ho7vCsgghSJQEcmy6uYpTgzd9czayOcxd89SH8
T55NpM+VFL/fvTc9YyZBz4wKdP8ZCzSyTCbcP8YvW1CzEWSYnWT4sVDa+vY7egQQ
9k/v50V4ECNq1D+3cythlN3V8KEzx0nRsI0gzjDDZ0fH162hCyiHjxIV6rzzuj+W
uJABHy+phSU3Lfw8WLg6/+8paUGiX6GoPGmprb8Tvypgvk7LFkycQhvZZFg+N9Xb
DmuK2sg6hiqrko3QWQQz1qUmuqA5l4ZZ9PUakkfZB2OGCdBSwborvhNIv7JzT78W
tHYury49BgLfbTVcLE7ozgQyD3D4imrhARF1fHcmDAfjSR70Rtx5HSRpWDjcq8Xi
SVr6r9jQATP6A3bWNhMN9jaje6/J5SQysgqV63o6fQgi0f0QdKdZETS6/x315SSe
eBcPw8eRiVzVX4853ZsPgUGv8P2QQqAA0/iMoZgpCTrk5YnHTnN/gzBGOkvQr5W5
MhYwOGAhRj8aKVayPAEK4MI7KwIhdzPt7VZ3Ok6Na/uLx1WDnQgKp62BiXMoQKA9
K7cqkfqngWL2nGs1d5NvxaFvkNJRruCAnelZmoC2kFuByZH8sI636JorG3DesR25
yJqc0YS560rSTc9ATcEO5hiybBZ07CuzpvgD/6AO0PysCySZaXAaw8Ouda7l93sP
wCSTv3iAOMeXL0wpzrw1IN0FpRgZPiP/lhV9NYhzEpJtGEYSSpsO3ChX1zsAmM7I
o72azqsHgRO68bZqLlN5symhU668BnUXIT4n5H7aRYAJhnVNo1IBLad9afDQ1hdA
IYDQ0YZo4xXATgmVtRFKSKkqR1wB0xWHpXFX+JsvI0HGqP3YCIDybOryhvlBYXUp
HYv/aMQ6pkSAPlrFm81fraSXW7ltJh5ExvFKMMstIus/jSU4+2kXVWbYECEzFaOs
oLmhMCyDxlx327jyS9Kkkj12dCTMp968NtilM/VD1PHTvMzY8VLrIdoj0yl81nCG
jkGk+6mWAQbdYytsC0WCKIdra9TpNq0xOnRK5bq9PIaL2QvcoB+eDWmFkTXrGyo4
HgoqoosfG4wbfhKQhPyPXfgMfVDCdMlMXr06O54jw5TJZAwGPXD8xzzL4nqUXb4I
ZlAqY6UvZs5Bvbt5jLStYMmjQsD1s/FdmZZyNYZgxbhVu8HX7xmhxKsMYARbiOCp
ITq02xqBepVBTTTZXMxqAeFxAOJPjSfeAlevNAai2LAMppr5k1boc3TW6Av9ATSH
vyQ7OjomBBQ619bzTU1Y1+sO18gRFY5xJU7/8Yy+v3oOnQVi58o1mZw3ILuX7aOX
fWtnwskoXmUxmx94Qz+CNdCgwrnyuKW9JihPzaqFSPx8zlXFa5IDpeDhmqbqLn1l
BGQllUJZ9Bm+FpZ9HUGOxA==
`protect END_PROTECTED
