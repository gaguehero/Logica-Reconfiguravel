`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BxeXpJlnrUqndqcHLo29p+i/s1gDHBNfY4kFfPFEWyXdpI7h7HYPjCGT3FF2c82F
mIUnc+7Ojgq474F1ThuSchNNDqvTJ4EAPxZ2hxs6jAnPCxRghQb2VEIZp0GDTV+v
wQ0+3XMPR9ds0Yc1yrQ4L5UV6DWu89lL5Gu7jx+R43haphxwYOhkB6RxOpNyWuMM
nShchFJItjpG/WlIXcir6Xly4uTSSyZyDvDJsG24rBE44JOmwTuhTDcHe/NCv9Ia
BuBg8qpV5s4SxcXoK3k2nfbnhpOlDhydep0jD/IQpUlregRvzgwG7KAtxRL8odAh
qSFSSUL8kBKBUoYHqomwiEG/K/aH7Vwoxn28/S/mgHWshuwqHn2N1IlBB9n2c/V3
lfXDHNgLJ193vozdYSDGuKbjJlBW6nMlrwu+C9SPE4UrsQMO0S34cTV2GXcYn2fN
YJTNxdAPcZayu0nGtmM5S7Aw4j/Po6us3T4xkesinW/0LvpQAbZOKIQqFTF+ppO7
0X5bV/Hwlo1GRfyyfao9e5L+nHgFlfcheaEa0SYMq6zcjPvyVJII3c+EtLLnsL0s
q8raC0CxhNYCNWOyz5AToi2aoIQ+LNOyCiph5fml22qYdLGu5bHROC76+Da7V8iE
SeMyGzVa2M7nDzH09oNZVg==
`protect END_PROTECTED
